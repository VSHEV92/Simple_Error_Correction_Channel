`include "Channel_Params.vh"

generate 
if (CHANNEL_PATTERN == 1) begin
     `define SYNDROME_TABLE_DEF SYNDROME_TABLE_7_4; 
end	
if (CHANNEL_PATTERN == 2) begin
	 `define SYNDROME_TABLE_DEF SYNDROME_TABLE_15_11; 
end	
if (CHANNEL_PATTERN == 3) begin
	 `define SYNDROME_TABLE_DEF SYNDROME_TABLE_15_7; 
end	
if (CHANNEL_PATTERN == 4) begin
	 `define SYNDROME_TABLE_DEF SYNDROME_TABLE_31_26; 
end
if (CHANNEL_PATTERN == 5) begin
	 `define SYNDROME_TABLE_DEF SYNDROME_TABLE_31_21; 
end
if (CHANNEL_PATTERN == 6) begin
	 `define SYNDROME_TABLE_DEF SYNDROME_TABLE_31_16; 
end			
endgenerate

parameter [0:`N_VAL*(2**(`N_VAL-`K_VAL))-1] SYNDROME_TABLE = `SYNDROME_TABLE_DEF;

parameter [0:7*(2**3)-1] SYNDROME_TABLE_7_4 = {
    7'b0000000,
    7'b0010000,
    7'b0100000,
    7'b0000001,
    7'b1000000,
    7'b0001000,
    7'b0000010,
    7'b0000100
};

parameter [0:15*(2**4)-1] SYNDROME_TABLE_15_11 = {
15'b000000000000000,
15'b000100000000000,
15'b001000000000000,
15'b000000000000001,
15'b010000000000000,
15'b000000000010000,
15'b000000000000010,
15'b000000001000000,
15'b100000000000000,
15'b000010000000000,
15'b000000000100000,
15'b000000000001000,
15'b000000000000100,
15'b000001000000000,
15'b000000010000000,
15'b000000100000000
};

parameter [0:15*(2**8)-1] SYNDROME_TABLE_15_7 = {
15'b000000000000000,
15'b000000010000000,
15'b000000100000000,
15'b000000110000000,
15'b000001000000000,
15'b000001010000000,
15'b000001100000000,
15'b000000000100010,
15'b000010000000000,
15'b000010010000000,
15'b000010100000000,
15'b000010110000000,
15'b000011000000000,
15'b000100000001000,
15'b000000001000100,
15'b000100100001000,
15'b000100000000000,
15'b000100010000000,
15'b000100100000000,
15'b011000000000010,
15'b000101000000000,
15'b000010000001000,
15'b000101100000000,
15'b001000000000101,
15'b000110000000000,
15'b000001000001000,
15'b001000000010000,
15'b100000001000010,
15'b000000010001000,
15'b000000000001000,
15'b001001000010000,
15'b000000100001000,
15'b001000000000000,
15'b001000010000000,
15'b001000100000000,
15'b010100000000010,
15'b001001000000000,
15'b100000000100001,
15'b110000000000100,
15'b000000000011000,
15'b001010000000000,
15'b010000000101000,
15'b000100000010000,
15'b000100010010000,
15'b001011000000000,
15'b001100000001000,
15'b010000000001010,
15'b000010000011000,
15'b001100000000000,
15'b010000100000010,
15'b000010000010000,
15'b010000000000010,
15'b010000000100000,
15'b010000010100000,
15'b010000100100000,
15'b000000000000101,
15'b000000100010000,
15'b000000001000001,
15'b000000000010000,
15'b000000010010000,
15'b010010000100000,
15'b001000000001000,
15'b000001000010000,
15'b001000100001000,
15'b010000000000000,
15'b010000010000000,
15'b010000100000000,
15'b010000110000000,
15'b010001000000000,
15'b010001010000000,
15'b101000000000100,
15'b010000000100010,
15'b010010000000000,
15'b000000000010010,
15'b010010100000000,
15'b000000100010010,
15'b100000000001001,
15'b010100000001000,
15'b000000000110000,
15'b000000010110000,
15'b010100000000000,
15'b100000000000001,
15'b100000001010000,
15'b001000000000010,
15'b001000000100000,
15'b100001000000001,
15'b001000100100000,
15'b001001000000010,
15'b010110000000000,
15'b100010000000001,
15'b011000000010000,
15'b001010000000010,
15'b100000000010100,
15'b010000000001000,
15'b000100000110000,
15'b010000100001000,
15'b011000000000000,
15'b011000010000000,
15'b100001000000100,
15'b000100000000010,
15'b000100000100000,
15'b000100010100000,
15'b100000000000100,
15'b100000010000100,
15'b100000001000000,
15'b000000000101000,
15'b100000101000000,
15'b100000000010001,
15'b100001001000000,
15'b000001000101000,
15'b000000000001010,
15'b000000010001010,
15'b000001000100000,
15'b000000100000010,
15'b000000010000010,
15'b000000000000010,
15'b000000000100000,
15'b000000010100000,
15'b000000100100000,
15'b000001000000010,
15'b100100001000000,
15'b010000001000001,
15'b010000000010000,
15'b000010000000010,
15'b000010000100000,
15'b011000000001000,
15'b010001000010000,
15'b000011000000010,
15'b100000000000000,
15'b100000010000000,
15'b100000100000000,
15'b100000110000000,
15'b100001000000000,
15'b100001010000000,
15'b100001100000000,
15'b100000000100010,
15'b100010000000000,
15'b100010010000000,
15'b100010100000000,
15'b000100001000010,
15'b100011000000000,
15'b100100000001000,
15'b100000001000100,
15'b000000000101100,
15'b100100000000000,
15'b010000000000001,
15'b000000000100100,
15'b010000100000001,
15'b100101000000000,
15'b000000000000110,
15'b000001000100100,
15'b000000100000110,
15'b100110000000000,
15'b100001000001000,
15'b101000000010000,
15'b000000001000010,
15'b000000001100000,
15'b100000000001000,
15'b000000101100000,
15'b100000100001000,
15'b101000000000000,
15'b101000010000000,
15'b000000000000011,
15'b000000010000011,
15'b101001000000000,
15'b000000000100001,
15'b010000000000100,
15'b100000000011000,
15'b010000001000000,
15'b010000011000000,
15'b100100000010000,
15'b010000000010001,
15'b010001001000000,
15'b000010000100001,
15'b010010000000100,
15'b000000000010110,
15'b101100000000000,
15'b011000000000001,
15'b100010000010000,
15'b110000000000010,
15'b110000000100000,
15'b010000001001000,
15'b010100000000100,
15'b100000000000101,
15'b100000100010000,
15'b100000001000001,
15'b100000000010000,
15'b100000010010000,
15'b001000001100000,
15'b101000000001000,
15'b100001000010000,
15'b000000000001011,
15'b110000000000000,
15'b000100000000001,
15'b110000100000000,
15'b000100100000001,
15'b110001000000000,
15'b000101000000001,
15'b001000000000100,
15'b001000010000100,
15'b001000001000000,
15'b100000000010010,
15'b001000101000000,
15'b001000000010001,
15'b000000000001001,
15'b000000010001001,
15'b100000000110000,
15'b000000001011000,
15'b000000010000001,
15'b000000000000001,
15'b000000001010000,
15'b000000100000001,
15'b101000000100000,
15'b000001000000001,
15'b001100000000100,
15'b000001100000001,
15'b001100001000000,
15'b000010000000001,
15'b000010001010000,
15'b010000001000010,
15'b000000000010100,
15'b110000000001000,
15'b000000100010100,
15'b000000001000101,
15'b000010001000000,
15'b001100000000001,
15'b000001000000100,
15'b100100000000010,
15'b000000100000100,
15'b010000000100001,
15'b000000000000100,
15'b000000010000100,
15'b000000001000000,
15'b000000011000000,
15'b000000101000000,
15'b000000000010001,
15'b000001001000000,
15'b000001011000000,
15'b000010000000100,
15'b000010010000100,
15'b100001000100000,
15'b001000000000001,
15'b100000010000010,
15'b100000000000010,
15'b100000000100000,
15'b000000001001000,
15'b000100000000100,
15'b100001000000010,
15'b000100001000000,
15'b001010000000001,
15'b110000000010000,
15'b000000000001100,
15'b100010000100000,
15'b000010001001000,
15'b000110000000100,
15'b000001000001100
};

parameter [0:31*(2**5)-1] SYNDROME_TABLE_31_26 = {
31'b0000000000000000000000000000000,
31'b0000100000000000000000000000000,
31'b0001000000000000000000000000000,
31'b0000000000000000010000000000000,
31'b0010000000000000000000000000000,
31'b0000000000000000000000000000001,
31'b0000000000000000100000000000000,
31'b0000000000000000000000001000000,
31'b0100000000000000000000000000000,
31'b0000001000000000000000000000000,
31'b0000000000000000000000000000010,
31'b0000000010000000000000000000000,
31'b0000000000000001000000000000000,
31'b0000000000000000000000000001000,
31'b0000000000000000000000010000000,
31'b0000000000001000000000000000000,
31'b1000000000000000000000000000000,
31'b0000000000000000000000000100000,
31'b0000010000000000000000000000000,
31'b0000000000000000001000000000000,
31'b0000000000000000000000000000100,
31'b0000000000000100000000000000000,
31'b0000000100000000000000000000000,
31'b0000000001000000000000000000000,
31'b0000000000000010000000000000000,
31'b0000000000100000000000000000000,
31'b0000000000000000000000000010000,
31'b0000000000000000000100000000000,
31'b0000000000000000000000100000000,
31'b0000000000000000000001000000000,
31'b0000000000010000000000000000000,
31'b0000000000000000000010000000000
};

parameter [0:31*(2**10)-1] SYNDROME_TABLE_31_21 = {
31'b0000000000000000000000000000000,
31'b0000000001000000000000000000000,
31'b0000000010000000000000000000000,
31'b0000000011000000000000000000000,
31'b0000000100000000000000000000000,
31'b0000000101000000000000000000000,
31'b0000000110000000000000000000000,
31'b0000100000000000100000000001000,
31'b0000001000000000000000000000000,
31'b0000001001000000000000000000000,
31'b0000001010000000000000000000000,
31'b1000000000000000000000000100100,
31'b0000001100000000000000000000000,
31'b0000000000000100000001000000000,
31'b0001000000000001000000000010000,
31'b0000000000000010000100000000000,
31'b0000010000000000000000000000000,
31'b0000010001000000000000000000000,
31'b0000010010000000000000000000000,
31'b0000000000000000001001000000000,
31'b0000010100000000000000000000000,
31'b1000000000010000000001000000000,
31'b1000000000100000100000000000000,
31'b1000000000001000000000001000000,
31'b0000011000000000000000000000000,
31'b0000000000000000100000000000010,
31'b0000000000001000000010000000000,
31'b0000100000010010000000000000000,
31'b0010000000000010000000000100000,
31'b1010000000000000000000010000000,
31'b0000000000000100001000000000000,
31'b0000000000000000000000000000101,
31'b0000100000000000000000000000000,
31'b0000100001000000000000000000000,
31'b0000100010000000000000000000000,
31'b1000000000000110000000000000000,
31'b0000100100000000000000000000000,
31'b0100000000000000000000100000100,
31'b0000000000000000010010000000000,
31'b0000000000000000100000000001000,
31'b0000101000000000000000000000000,
31'b0100000000100000000000010000000,
31'b0010000000000000001000000000100,
31'b1000000000000000010000001000000,
31'b1000000000000100000100000000000,
31'b0000000000000001000000000000001,
31'b1000000000000010000001000000000,
31'b0000100000000010000100000000000,
31'b0000110000000000000000000000000,
31'b1000000000100000000000000001000,
31'b0000000000000001000000000000100,
31'b0000100000000000001001000000000,
31'b0000000000010000000100000000000,
31'b0100000000000000000001001000000,
31'b0001000000100100000000000000000,
31'b0100000000011000000000000000000,
31'b0100000000000100000000001000000,
31'b1000000000000001000000000100000,
31'b0100000000000000000000100000001,
31'b0000000000010010000000000000000,
31'b0000000000001000010000000000000,
31'b1000000000000010001000000000000,
31'b0000000000000000000000000001010,
31'b0100000000000000010100000000000,
31'b0001000000000000000000000000000,
31'b0001000001000000000000000000000,
31'b0001000010000000000000000000000,
31'b0000000000000010100000000000000,
31'b0001000100000000000000000000000,
31'b0010000000000000000001000010000,
31'b0010000000000000000000000100010,
31'b1000000000000100000000000001000,
31'b0001001000000000000000000000000,
31'b0001001001000000000000000000000,
31'b1000000000000000000001000001000,
31'b0000100000000000000100000001000,
31'b0000000000000000100100000000000,
31'b0010100000001000000000000000000,
31'b0000000000000001000000000010000,
31'b0100000000001000100000000000000,
31'b0001010000000000000000000000000,
31'b0010000000000000010000000000000,
31'b1000000001000000000000100000000,
31'b1000000000000000000000100000000,
31'b0100000000000000010000000001000,
31'b0000000000000000000100000000010,
31'b0100000000001000000000000000010,
31'b1000000100000000000000100000000,
31'b0001011000000000000000000000000,
31'b1000000000000000001000000001000,
31'b0000000000000010000000000000010,
31'b1000001000000000000000100000000,
31'b0000100000000000000000000010100,
31'b0100100000000000000000000100000,
31'b0001000000000100001000000000000,
31'b0000000000010000000000000001000,
31'b0001100000000000000000000000000,
31'b0000000000010000000000000000010,
31'b0001100010000000000000000000000,
31'b0000000000000000000000000010001,
31'b0000000000000010000000000001000,
31'b0010001000001000000000000000000,
31'b0001000000000000010010000000000,
31'b0000000000000000000000011000000,
31'b0000000000100000001000000000000,
31'b1100000000000000000000000000001,
31'b1000000000000000000010010000000,
31'b0000000000000000000100000001000,
31'b0010000001001000000000000000000,
31'b0010000000001000000000000000000,
31'b1000000000110000000000000000000,
31'b0010000010001000000000000000000,
31'b1000000000001000000000010000000,
31'b0010100000000000010000000000000,
31'b0100000000000000000010000001000,
31'b1000100000000000000000100000000,
31'b1000000000000000000001000000010,
31'b0100001000000000000000000100000,
31'b0000000000100100000000000000000,
31'b0010000000000000000010000000000,
31'b0000000000010000100000000000000,
31'b1000000000000100000000000000010,
31'b1010000000000000000000001000000,
31'b0000000000100000000001000000000,
31'b0000000000000000000000000010100,
31'b0100000000000000000000000100000,
31'b1000000000000000101000000000000,
31'b0100000010000000000000000100000,
31'b0010000000000000000000000000000,
31'b0010000001000000000000000000000,
31'b0010000010000000000000000000000,
31'b0010000011000000000000000000000,
31'b0010000100000000000000000000000,
31'b0100000000000000000000000001000,
31'b0000000000000101000000000000000,
31'b1000000000000000000100000000001,
31'b0010001000000000000000000000000,
31'b0010001001000000000000000000000,
31'b0100000000000000000010000100000,
31'b0000000000000001000001000000000,
31'b0100000000000000000000001000100,
31'b1000010000000000000000010000000,
31'b0001000000000000000000110000000,
31'b1000000000000000000000000011000,
31'b0010010000000000000000000000000,
31'b0001000000000000010000000000000,
31'b0010010010000000000000000000000,
31'b0000000000000000000100000100000,
31'b0010010100000000000000000000000,
31'b1000001000000000000000010000000,
31'b0001000000000000001000000010000,
31'b1000000000000010000000000000100,
31'b0000000000000001001000000000000,
31'b1000000100000000000000010000000,
31'b0101000000010000000000000000000,
31'b0100100000000000000000000000010,
31'b0000000000000010000000000100000,
31'b1000000000000000000000010000000,
31'b1000000000010001000000000000000,
31'b1000000010000000000000010000000,
31'b0010100000000000000000000000000,
31'b1000000000000000001000000100000,
31'b0100000000000000100000000000000,
31'b0100000001000000100000000000000,
31'b1000000000000000000010100000000,
31'b1000000000000011000000000000000,
31'b0000000000000000000001000000001,
31'b0000000000010000000000000100000,
31'b1000000000000000100000000010000,
31'b0000000000000000000000101000000,
31'b0000000000000000001000000000100,
31'b0000000000000100000000000000001,
31'b1000000000010000000000000000100,
31'b0001000000001000000000000000000,
31'b0101000000000000000100000000000,
31'b0001000010001000000000000000000,
31'b0010110000000000000000000000000,
31'b1000000000000000000000000010010,
31'b1000000000000000000001000100000,
31'b1000000000010000000000000000001,
31'b0000000000000100000000000000100,
31'b0000000000000000001000000000001,
31'b0001000001000000000010000000000,
31'b0001000000000000000010000000000,
31'b0001000000000000000000000101000,
31'b0000000000000000000001000000100,
31'b1001000000000000000000001000000,
31'b0100000000000000000000000000010,
31'b0010000000001000010000000000000,
31'b1000100000000000000000010000000,
31'b0000000000100000000000000010000,
31'b1000000000000100000000000100000,
31'b0011000000000000000000000000000,
31'b0000010000000000010000000000000,
31'b0000000000100000000000000000100,
31'b0010000000000010100000000000000,
31'b0011000100000000000000000000000,
31'b0000000000000000000001000010000,
31'b0000000000000000000000000100010,
31'b0000110000000000000010000000000,
31'b0000000000000100000000000010000,
31'b1000000000100000000000000100000,
31'b0100010000010000000000000000000,
31'b1000000000000000100000000000001,
31'b0010000000000000100100000000000,
31'b0000100000001000000000000000000,
31'b0000000000000000000000110000000,
31'b1100000000000000000001000000000,
31'b0000000001000000010000000000000,
31'b0000000000000000010000000000000,
31'b1000000000000000000000000000011,
31'b0000000010000000010000000000000,
31'b1000000000000000100000000000100,
31'b0000000100000000010000000000000,
31'b0000000000000000001000000010000,
31'b0000100000000000000010000000000,
31'b0100000010010000000000000000000,
31'b0000001000000000010000000000000,
31'b0100000000010000000000000000000,
31'b0100000001010000000000000000000,
31'b1100000000000000001000000000000,
31'b0000000000100000000000000000001,
31'b0100000100010000000000000000000,
31'b0000000000000000100000000100000,
31'b0100000001000010000000000000000,
31'b0100000000000010000000000000000,
31'b0101000000000000100000000000000,
31'b0100000010000010000000000000000,
31'b1000000000000000000100000010000,
31'b0000001000001000000000000000000,
31'b1000000000000001100000000000000,
31'b0000010000000000000010000000000,
31'b0010000000100000001000000000000,
31'b0000000100001000000000000000000,
31'b1000010000000000000000001000000,
31'b1000000000000010000000000010000,
31'b0000000001001000000000000000000,
31'b0000000000001000000000000000000,
31'b0100000000000000000100000000000,
31'b0000000010001000000000000000000,
31'b0000000000100001000000000000000,
31'b0000100000000000010000000000000,
31'b1000001000000000000000001000000,
31'b0000000100000000000010000000000,
31'b0100000000000000000000010000001,
31'b0000000010000000000010000000000,
31'b0000000001000000000010000000000,
31'b0000000000000000000010000000000,
31'b0000000000000000000000000101000,
31'b0001000000000000000001000000100,
31'b1000000000000000000000001000000,
31'b1000000001000000000000001000000,
31'b0010000000000000000000000010100,
31'b0000010000001000000000000000000,
31'b1000000100000000000000001000000,
31'b0000001000000000000010000000000,
31'b0100000000000000000000000000000,
31'b0100000001000000000000000000000,
31'b0100000010000000000000000000000,
31'b0000000000001000000100000000000,
31'b0100000100000000000000000000000,
31'b0010000000000000000000000001000,
31'b0100000110000000000000000000000,
31'b0010000010000000000000000001000,
31'b0100001000000000000000000000000,
31'b0100001001000000000000000000000,
31'b1000000000000000000000000010000,
31'b0000000000010000010000000000000,
31'b0000000000001010000000000000000,
31'b1000000000000000011000000000000,
31'b1000000100000000000000000010000,
31'b0100000000000010000100000000000,
31'b0100010000000000000000000000000,
31'b0100010001000000000000000000000,
31'b0100010010000000000000000000000,
31'b1000000000000100010000000000000,
31'b1000000000000000000100001000000,
31'b0010010000000000000000000001000,
31'b0000000000000010000010000000000,
31'b0000000000000001000000100000000,
31'b1000000000000000000000010001000,
31'b0000000000000000000110000000000,
31'b1000010000000000000000000010000,
31'b1000000000000010000000001000000,
31'b0010000000000000000001100000000,
31'b0001100000000000000000000100000,
31'b1000000000000000010001000000000,
31'b0100000000000000000000000000101,
31'b0100100000000000000000000000000,
31'b0100100001000000000000000000000,
31'b0010000000000000100000000000000,
31'b0010000001000000100000000000000,
31'b0100100100000000000000000000000,
31'b0000000000000000000000100000100,
31'b0000000000000000001000001000000,
31'b0100000000000000100000000001000,
31'b0100101000000000000000000000000,
31'b0000000000100000000000010000000,
31'b1000100000000000000000000010000,
31'b1000000000000000001010000000000,
31'b0010000000000000010000000100000,
31'b0000000000010000000010000000000,
31'b1000000000000000000000100100000,
31'b1000000000001100000000000000000,
31'b0000000000000010010000000000000,
31'b1000000000001000001000000000000,
31'b0100000000000001000000000000100,
31'b0010001000000000000000000000010,
31'b1010000000100000000000000000000,
31'b0000000000000000000001001000000,
31'b1001000000000000000000000000100,
31'b0000000000011000000000000000000,
31'b0000000000000100000000001000000,
31'b0010000010000000000000000000010,
31'b0000000000000000000000100000001,
31'b0010000000000000000000000000010,
31'b0100000000001000010000000000000,
31'b0001000000000000000000000100000,
31'b0100000000000000000000000001010,
31'b0000000000000000010100000000000,
31'b0101000000000000000000000000000,
31'b0000000000000000001000010000000,
31'b1010000000000100000000000000000,
31'b1000000000100000000010000000000,
31'b1000000000000001000000000000000,
31'b1000000001000001000000000000000,
31'b1000000010000001000000000000000,
31'b1000000000010000000000010000000,
31'b0101001000000000000000000000000,
31'b1000100000000000000000000000001,
31'b1001000000000000000000000010000,
31'b0001000000010000010000000000000,
31'b0000000000000000000010000000010,
31'b0000110000000000000000000100000,
31'b0000000000100000000000001000000,
31'b0000000000001000100000000000000,
31'b0101010000000000000000000000000,
31'b0110000000000000010000000000000,
31'b0000000000000000000001010000000,
31'b1100000000000000000000100000000,
31'b0000000000000000010000000001000,
31'b0000000000000000100010000000000,
31'b0000000000001000000000000000010,
31'b0001000000000001000000100000000,
31'b1000000000000000100000001000000,
31'b0000000000000000000000100010000,
31'b0010000000010000000000000000000,
31'b0010000001010000000000000000000,
31'b1010000000000000001000000000000,
31'b0000100000000000000000000100000,
31'b0010000100010000000000000000000,
31'b0000000000000100000000010000000,
31'b0101100000000000000000000000000,
31'b0010000000000010000000000000000,
31'b0011000000000000100000000000000,
31'b0100000000000000000000000010001,
31'b1000100000000001000000000000000,
31'b1000000000100000010000000000000,
31'b1000010000000000000000000000100,
31'b0100000000000000000000011000000,
31'b0000000000001000000000000001000,
31'b1000000000000000000000000000001,
31'b0000000000000000010000000000010,
31'b1000000010000000000000000000001,
31'b0010000010000000000100000000000,
31'b0000010000000000000000000100000,
31'b0010000000000000000100000000000,
31'b0010000001000000000100000000000,
31'b0010000000000000000000001010000,
31'b0010010000000010000000000000000,
31'b0000000000000000000010000001000,
31'b0000000000000000110000000000000,
31'b1000000010000000000000000000100,
31'b0000001000000000000000000100000,
31'b1000000000000000000000000000100,
31'b1000000001000000000000000000100,
31'b0100000000010000100000000000000,
31'b0000000100000000000000000100000,
31'b0010100000010000000000000000000,
31'b0100000000100000000001000000000,
31'b0000000001000000000000000100000,
31'b0000000000000000000000000100000,
31'b1000001000000000000000000000100,
31'b0000000010000000000000000100000,
31'b0110000000000000000000000000000,
31'b0000000100000000000000000001000,
31'b0000100000000000100000000000000,
31'b0010000000001000000100000000000,
31'b0000000001000000000000000001000,
31'b0000000000000000000000000001000,
31'b0100000000000101000000000000000,
31'b0000000010000000000000000001000,
31'b0110001000000000000000000000000,
31'b1000000000010000000000100000000,
31'b0000000000000000000010000100000,
31'b0100000000000001000001000000000,
31'b0000000000000000000000001000100,
31'b0000001000000000000000000001000,
31'b0001100000000000000100000000000,
31'b0000000000000000001000100000000,
31'b0000000000001000000000000100000,
31'b0000000000000100000000100000000,
31'b0001001000010000000000000000000,
31'b0000000000000000000000001000001,
31'b1000100000100000000000000000000,
31'b0000010000000000000000000001000,
31'b0010000000000010000010000000000,
31'b0000000000000000000000010010000,
31'b0100000000000001001000000000000,
31'b0010000000000000000110000000000,
31'b0001000000010000000000000000000,
31'b0000100000000000000000000000010,
31'b0000000000000000000001100000000,
31'b1100000000000000000000010000000,
31'b1000000000000000000010000000001,
31'b0000100100000000000000000000010,
31'b0000000010000000100000000000000,
31'b0001000000000010000000000000000,
31'b0000000000000000100000000000000,
31'b0000000001000000100000000000000,
31'b1000010000100000000000000000000,
31'b0000100000000000000000000001000,
31'b0000000100000000100000000000000,
31'b1000000000000000010000000000100,
31'b0000001010000000100000000000000,
31'b1000000000001001000000000000000,
31'b0000001000000000100000000000000,
31'b0000010000000000000000000000010,
31'b0000000000000000010000000100000,
31'b0101000000001000000000000000000,
31'b0001000000000000000100000000000,
31'b0001000001000000000100000000000,
31'b1000000100100000000000000000000,
31'b0001010000000010000000000000000,
31'b0000010000000000100000000000000,
31'b0000001000000000000000000000010,
31'b1000000000100000000000000000000,
31'b1000000001100000000000000000000,
31'b1000000010100000000000000000000,
31'b0101000000000000000010000000000,
31'b1000000000000000010000000000001,
31'b0000000010000000000000000000010,
31'b0000000001000000000000000000010,
31'b0000000000000000000000000000010,
31'b1000001000100000000000000000000,
31'b1000000000000000000100100000000,
31'b0000000000000001000000001000000,
31'b0000000100000000000000000000010,
31'b1000000010000100000000000000000,
31'b0000100000000010000000000000000,
31'b1000000000000100000000000000000,
31'b1000000001000100000000000000000,
31'b1010000000000001000000000000000,
31'b0001000000000000000000000001000,
31'b1000000100000100000000000000000,
31'b1000001000000000000001000000000,
31'b0100000000000100000000000010000,
31'b0000101000000010000000000000000,
31'b0000010000010000000000000000000,
31'b1000000100000000000001000000000,
31'b1000010000000000001000000000000,
31'b1000000010000000000001000000000,
31'b0000100000000000000100000000000,
31'b1000000000000000000001000000000,
31'b0100000001000000010000000000000,
31'b0100000000000000010000000000000,
31'b0000001000010000000000000000000,
31'b0100000010000000010000000000000,
31'b1000001000000000001000000000000,
31'b0100000100000000010000000000000,
31'b1000000000000000000000100001000,
31'b0100100000000000000010000000000,
31'b0000000010010000000000000000000,
31'b0000000000000001000000010000000,
31'b0000000000010000000000000000000,
31'b0000000001010000000000000000000,
31'b1000000000000000001000000000000,
31'b1000000001000000001000000000000,
31'b0000000100010000000000000000000,
31'b1000010000000000000001000000000,
31'b0000000001000010000000000000000,
31'b0000000000000010000000000000000,
31'b0001000000000000100000000000000,
31'b0000000010000010000000000000000,
31'b0000010000000000000000010000001,
31'b0000000100000010000000000000000,
31'b0000001000000000000100000000000,
31'b0000000000100000000000100000000,
31'b1000000000000000000000100000010,
31'b0000001000000010000000000000000,
31'b0000000100000000000100000000000,
31'b0000000000000000000000010000100,
31'b0000000010000000000100000000000,
31'b0100000000001000000000000000000,
31'b0000000000000000000100000000000,
31'b0000000001000000000100000000000,
31'b0000000000000000000000001010000,
31'b0000010000000010000000000000000,
31'b0010000000000000000010000001000,
31'b0100000100000000000010000000000,
31'b0000000000000000000000010000001,
31'b0100000010000000000010000000000,
31'b1010000000000000000000000000100,
31'b0100000000000000000010000000000,
31'b0100000000000000000000000101000,
31'b0010000100000000000000000100000,
31'b0000100000010000000000000000000,
31'b0001000000000000000000000000010,
31'b1000100000000000001000000000000,
31'b0010000000000000000000000100000,
31'b0000010000000000000100000000000,
31'b0100001000000000000010000000000,
31'b1000000000000000000000000000000,
31'b1000000001000000000000000000000,
31'b1000000010000000000000000000000,
31'b1000000011000000000000000000000,
31'b1000000100000000000000000000000,
31'b1000000101000000000000000000000,
31'b0000000000010000001000000000000,
31'b0010000000000000000100000000001,
31'b1000001000000000000000000000000,
31'b1000001001000000000000000000000,
31'b0100000000000000000000000010000,
31'b0000000000000000000000000100100,
31'b1000001100000000000000000000000,
31'b0000000000000000000010001000000,
31'b0100000100000000000000000010000,
31'b0000000000100000000000000000010,
31'b1000010000000000000000000000000,
31'b1000010001000000000000000000000,
31'b1000010010000000000000000000000,
31'b0001000000000000000000100000000,
31'b0000000000000000000000000100001,
31'b0000000000010000000001000000000,
31'b0000000000100000100000000000000,
31'b0000000000001000000000001000000,
31'b0000000000010100000000000000000,
31'b1000000000000000100000000000010,
31'b1000000000001000000010000000000,
31'b0100000000000010000000001000000,
31'b0010000001000000000000010000000,
31'b0010000000000000000000010000000,
31'b1000000000000100001000000000000,
31'b1000000000000000000000000000101,
31'b1000100000000000000000000000000,
31'b0000000000000000000101000000000,
31'b1000100010000000000000000000000,
31'b0000000000000110000000000000000,
31'b1000100100000000000000000000000,
31'b0010000000000011000000000000000,
31'b1000000000000000010010000000000,
31'b1000000000000000100000000001000,
31'b1000101000000000000000000000000,
31'b0101000000000000000000000000001,
31'b0100100000000000000000000010000,
31'b0000000000000000010000001000000,
31'b0000000000000100000100000000000,
31'b1000000000000001000000000000001,
31'b0000000000000010000001000000000,
31'b0100000000001100000000000000000,
31'b1000110000000000000000000000000,
31'b0000000000100000000000000001000,
31'b0000000000000000001100000000000,
31'b0010000000010000000000000000001,
31'b1000000000010000000100000000000,
31'b0100000000000100000010000000000,
31'b0101000000000000000000000000100,
31'b0001000000000000000000000110000,
31'b0100000000000000000011000000000,
31'b0000000000000001000000000100000,
31'b0011000000000000000000001000000,
31'b1000000000010010000000000000000,
31'b1000000000001000010000000000000,
31'b0000000000000010001000000000000,
31'b1000000000000000000000000001010,
31'b0100000000000000100000010000000,
31'b1001000000000000000000000000000,
31'b1001000001000000000000000000000,
31'b1001000010000000000000000000000,
31'b0000010000000000000000100000000,
31'b0100000000000001000000000000000,
31'b0100000001000001000000000000000,
31'b0100000010000001000000000000000,
31'b0000000000000100000000000001000,
31'b1001001000000000000000000000000,
31'b0100100000000000000000000000001,
31'b0000000000000000000001000001000,
31'b0010000000000000100000000000001,
31'b0000000000000000010000010000000,
31'b0010000000000000000000000000110,
31'b1000000000000001000000000010000,
31'b0110000000000000000001000000000,
31'b1001010000000000000000000000000,
31'b0000000010000000000000100000000,
31'b0000000001000000000000100000000,
31'b0000000000000000000000100000000,
31'b0100010000000001000000000000000,
31'b0000000000100010000000000000000,
31'b0100100000000000000000000000100,
31'b0000000100000000000000100000000,
31'b0100000000000000100000001000000,
31'b0000000000000000001000000001000,
31'b0000000000100000000100000000000,
31'b0000001000000000000000100000000,
31'b0110000000000000001000000000000,
31'b0011000000000000000000010000000,
31'b0000100000000000101000000000000,
31'b1000000000010000000000000001000,
31'b0000000000000100100000000000000,
31'b1000000000010000000000000000010,
31'b0000001000000000000010010000000,
31'b1000000000000000000000000010001,
31'b1000000000000010000000000001000,
31'b0100000000100000010000000000000,
31'b0100010000000000000000000000100,
31'b0000000000000000001000000000010,
31'b1000000000100000001000000000000,
31'b0100000000000000000000000000001,
31'b0000000000000000000010010000000,
31'b1000000000000000000100000001000,
31'b0010000000000000000000000001001,
31'b0000000000000000100001000000000,
31'b0000000000110000000000000000000,
31'b0000001000000000001000000000010,
31'b0000000000001000000000010000000,
31'b0001000000100000000000000001000,
31'b0100000100000000000000000000100,
31'b0000100000000000000000100000000,
31'b0000000000000000000001000000010,
31'b0000100000100010000000000000000,
31'b0100000000000000000000000000100,
31'b0000000000000000000000000110000,
31'b1000000000010000100000000000000,
31'b0000000000000100000000000000010,
31'b0010000000000000000000001000000,
31'b1000000000100000000001000000000,
31'b1000000000000000000000000010100,
31'b1100000000000000000000000100000,
31'b0000000000000000101000000000000,
31'b0100000000000000000000001001000,
31'b1010000000000000000000000000000,
31'b1010000001000000000000000000000,
31'b0000000000000000010000100000000,
31'b0000000100000000000100000000001,
31'b1010000100000000000000000000000,
31'b1100000000000000000000000001000,
31'b1000000000000101000000000000000,
31'b0000000000000000000100000000001,
31'b0000000000000010000000000000001,
31'b0100000000010000000000100000000,
31'b0110000000000000000000000010000,
31'b1000000000000001000001000000000,
31'b0000100000010000000000000000100,
31'b0000010000000000000000010000000,
31'b0000010000010001000000000000000,
31'b0000000000000000000000000011000,
31'b1010010000000000000000000000000,
31'b1001000000000000010000000000000,
31'b0001000000000000000000000000011,
31'b1000000000000000000100000100000,
31'b0100100000100000000000000000000,
31'b0000001000000000000000010000000,
31'b0010000000100000100000000000000,
31'b0000000000000010000000000000100,
31'b0000000000000000000100000000100,
31'b0000000100000000000000010000000,
31'b0001100000000000000000001000000,
31'b0100000000001000000000000000100,
31'b0000000001000000000000010000000,
31'b0000000000000000000000010000000,
31'b0000000000010001000000000000000,
31'b0000000010000000000000010000000,
31'b1010100000000000000000000000000,
31'b0000000000000000001000000100000,
31'b1100000000000000100000000000000,
31'b0010000000000110000000000000000,
31'b0000000000000000000010100000000,
31'b0000000000000011000000000000000,
31'b1000000000000000000001000000001,
31'b1000000000010000000000000100000,
31'b0000000000000000100000000010000,
31'b1000000000000000000000101000000,
31'b0000000000000001000100000000000,
31'b1000000000000100000000000000001,
31'b0000000000010000000000000000100,
31'b1001000000001000000000000000000,
31'b0010000000000010000001000000000,
31'b0000100000000000000000000011000,
31'b0100000100100000000000000000000,
31'b0000000000000000000000000010010,
31'b0000000000000000000001000100000,
31'b0000000000010000000000000000001,
31'b0100000000100000000000000000000,
31'b1000000000000000001000000000001,
31'b0100000010100000000000000000000,
31'b1001000000000000000010000000000,
31'b0100000000000000010000000000001,
31'b1000000000000000000001000000100,
31'b0001000000000000000000001000000,
31'b1100000000000000000000000000010,
31'b0100001000100000000000000000000,
31'b0000100000000000000000010000000,
31'b0000000000001000000000100000000,
31'b0000000000000100000000000100000,
31'b1011000000000000000000000000000,
31'b0000000000000001000000000001000,
31'b0100000000000100000000000000000,
31'b0100000001000100000000000000000,
31'b0110000000000001000000000000000,
31'b1000000000000000000001000010000,
31'b1000000000000000000000000100010,
31'b0100001000000000000001000000000,
31'b1000000000000100000000000010000,
31'b0000000000100000000000000100000,
31'b0100001000000100000000000000000,
31'b0000000000000000100000000000001,
31'b0100010000000000001000000000000,
31'b0000000000000000000000000000110,
31'b1000000000000000000000110000000,
31'b0100000000000000000001000000000,
31'b0000000000010000000000000010000,
31'b1000000000000000010000000000000,
31'b0000000000000000000000000000011,
31'b0010000000000000000000100000000,
31'b0000000000000000100000000000100,
31'b1000000100000000010000000000000,
31'b1000000000000000001000000010000,
31'b1000100000000000000010000000000,
31'b0100000100000000001000000000000,
31'b1000001000000000010000000000000,
31'b0000100000000000000000001000000,
31'b0100000000000000010000000010000,
31'b0100000000000000001000000000000,
31'b0001000000000000000000010000000,
31'b0100000010000000001000000000000,
31'b1000000000000000100000000100000,
31'b0100000000000000000000010100000,
31'b1100000000000010000000000000000,
31'b0100100000000100000000000000000,
31'b0000010000000000000000000001100,
31'b0000000000000000000100000010000,
31'b1000001000001000000000000000000,
31'b0000000000000001100000000000000,
31'b1000010000000000000010000000000,
31'b0100000000000000000000100000010,
31'b1000000100001000000000000000000,
31'b0000010000000000000000001000000,
31'b0000000000000010000000000010000,
31'b0000000000000000000000000001001,
31'b1000000000001000000000000000000,
31'b1100000000000000000100000000000,
31'b1000000010001000000000000000000,
31'b1000000000100001000000000000000,
31'b1000100000000000010000000000000,
31'b0000001000000000000000001000000,
31'b0000000000000000000000000001100,
31'b0101000000100000000000000000000,
31'b1000000010000000000010000000000,
31'b1000000001000000000010000000000,
31'b1000000000000000000010000000000,
31'b0000000010000000000000001000000,
31'b0010000000000100000000000000010,
31'b0000000000000000000000001000000,
31'b0000000001000000000000001000000,
31'b0100100000000000001000000000000,
31'b1000010000001000000000000000000,
31'b0000000100000000000000001000000,
31'b0000000000000001000000000000010,
31'b1100000000000000000000000000000,
31'b1100000001000000000000000000000,
31'b0000001000000000000000000010000,
31'b1000000000001000000100000000000,
31'b0001000000000001000000000000000,
31'b1010000000000000000000000001000,
31'b0100000000010000001000000000000,
31'b0010000000000000000000001100000,
31'b0000000010000000000000000010000,
31'b0010000000010000000000100000000,
31'b0000000000000000000000000010000,
31'b0000000001000000000000000010000,
31'b1000000000001010000000000000000,
31'b0000000000000000011000000000000,
31'b0000000100000000000000000010000,
31'b0100000000100000000000000000010,
31'b1100010000000000000000000000000,
31'b0000100000001000001000000000000,
31'b0000011000000000000000000010000,
31'b0000000000000100010000000000000,
31'b0000000000000000000100001000000,
31'b0100000000010000000001000000000,
31'b1000000000000010000010000000000,
31'b1000000000000001000000100000000,
31'b0000000000000000000000010001000,
31'b1000000000000000000110000000000,
31'b0000010000000000000000000010000,
31'b0000000000000010000000001000000,
31'b0011000000000000001000000000000,
31'b0110000000000000000000010000000,
31'b0000000000000000010001000000000,
31'b0000100000000000100000010000000,
31'b0000000000010000000000001000000,
31'b0100000000000000000101000000000,
31'b0000000000001000000001000000000,
31'b0100000000000110000000000000000,
31'b0010010000100000000000000000000,
31'b1000000000000000000000100000100,
31'b0000000000000000000000010000010,
31'b0010000000000000010000000000100,
31'b0001000001000000000000000000001,
31'b0001000000000000000000000000001,
31'b0000100000000000000000000010000,
31'b0000000000000000001010000000000,
31'b0100000000000100000100000000000,
31'b1000000000010000000010000000000,
31'b0000000000000000000000100100000,
31'b0000000000001100000000000000000,
31'b1000000000000010010000000000000,
31'b0000000000001000001000000000000,
31'b0100000000000000001100000000000,
31'b0010000000000001000010000000000,
31'b0010000000100000000000000000000,
31'b0000000000000100000010000000000,
31'b0001000000000000000000000000100,
31'b1000000000011000000000000000000,
31'b0000000000000000000011000000000,
31'b0100000000000001000000000100000,
31'b1000000000000000000000100000001,
31'b1010000000000000000000000000010,
31'b0010001000100000000000000000000,
31'b1001000000000000000000000100000,
31'b0001001000000000000000000000100,
31'b0000000000000000100000010000000,
31'b0000000100000001000000000000000,
31'b0000000000000000000000001000010,
31'b0010000000000100000000000000000,
31'b0000000000100000000010000000000,
31'b0000000000000001000000000000000,
31'b0000000001000001000000000000000,
31'b0000000010000001000000000000000,
31'b0000000000010000000000010000000,
31'b0001000010000000000000000010000,
31'b0000100000000000000000000000001,
31'b0001000000000000000000000010000,
31'b0010000100000000000001000000000,
31'b0000001000000001000000000000000,
31'b0010000010000000000001000000000,
31'b1000000000100000000000001000000,
31'b0010000000000000000001000000000,
31'b0000010100000001000000000000000,
31'b0100000010000000000000100000000,
31'b1000000000000000000001010000000,
31'b0100000000000000000000100000000,
31'b0000010000000001000000000000000,
31'b1000000000000000100010000000000,
31'b0000100000000000000000000000100,
31'b0100000100000000000000100000000,
31'b0000000000000000100000001000000,
31'b0000000000101000000000000000000,
31'b1010000000010000000000000000000,
31'b0100001000000000000000100000000,
31'b0010000000000000001000000000000,
31'b1000100000000000000000000100000,
31'b0010000010000000001000000000000,
31'b1000000000000100000000010000000,
31'b0100000000000100100000000000000,
31'b0000001000000000000000000000001,
31'b0010100000000100000000000000000,
31'b0000100000100000000010000000000,
31'b0000100000000001000000000000000,
31'b0000000000100000010000000000000,
31'b0000010000000000000000000000100,
31'b0100000000000000001000000000010,
31'b0000000001000000000000000000001,
31'b0000000000000000000000000000001,
31'b1000000000000000010000000000010,
31'b0000000010000000000000000000001,
31'b0000101000000001000000000000000,
31'b0000000100000000000000000000001,
31'b1010000000000000000100000000000,
31'b0010100000000000000001000000000,
31'b0100000000001000000000010000000,
31'b0010000000000000100000100000000,
31'b0000000100000000000000000000100,
31'b0000000000000000000100010000000,
31'b0000000010000000000000000000100,
31'b1000001000000000000000000100000,
31'b0000000000000000000000000000100,
31'b0000000001000000000000000000100,
31'b0001000000000000000011000000000,
31'b0000010000000000000000000000001,
31'b0110000000000000000000001000000,
31'b0000010010000000000000000000001,
31'b0000000000000010000000010000000,
31'b1000000000000000000000000100000,
31'b0000001000000000000000000000100,
31'b0000000000000000000000001001000,
31'b1110000000000000000000000000000,
31'b0000000000000000000010000000100,
31'b0001000000000100000000000000000,
31'b0001000001000100000000000000000,
31'b0000000000001000000000000000001,
31'b1000000000000000000000000001000,
31'b0001000100000100000000000000000,
31'b0000000000000000000000001100000,
31'b0100000000000010000000000000001,
31'b0000000000010000000000100000000,
31'b0010000000000000000000000010000,
31'b0010000001000000000000000010000,
31'b1000000000000000000000001000100,
31'b1000001000000000000000000001000,
31'b0010000100000000000000000010000,
31'b0001000000000000000001000000000,
31'b1000000000001000000000000100000,
31'b1000000000000100000000100000000,
31'b0001010000000100000000000000000,
31'b1000000000000000000000001000001,
31'b0000100000100000000000000000000,
31'b0000000000000001010000000000000,
31'b0001000000000000000000100001000,
31'b1000000000000000000000010010000,
31'b0100000000000000000100000000100,
31'b0100000100000000000000010000000,
31'b1001000000010000000000000000000,
31'b0000000000001000000000000000100,
31'b0001000000000000001000000000000,
31'b0100000000000000000000010000000,
31'b0000000000000000000010000000001,
31'b0100000010000000000000010000000,
31'b1000000010000000100000000000000,
31'b1001000000000010000000000000000,
31'b1000000000000000100000000000000,
31'b1000000001000000100000000000000,
31'b0000010000100000000000000000000,
31'b1000100000000000000000000001000,
31'b1000000100000000100000000000000,
31'b0000000000000000010000000000100,
31'b0100000000000000100000000010000,
31'b0000000000001001000000000000000,
31'b1000001000000000100000000000000,
31'b1000010000000000000000000000010,
31'b1000000000000000010000000100000,
31'b0000010000000000000100100000000,
31'b1001000000000000000100000000000,
31'b0010000000001100000000000000000,
31'b0000000100100000000000000000000,
31'b0100000000000000000000000010010,
31'b0000000000000010000000100000000,
31'b0000000000000001000010000000000,
31'b0000000000100000000000000000000,
31'b0000000001100000000000000000000,
31'b0000000010100000000000000000000,
31'b0000010000000000010000000000100,
31'b0000000000000000010000000000001,
31'b1000000010000000000000000000010,
31'b1000000001000000000000000000010,
31'b1000000000000000000000000000010,
31'b0000001000100000000000000000000,
31'b0000000000000000000100100000000,
31'b1000000000000001000000001000000,
31'b1000000100000000000000000000010,
31'b0000000010000100000000000000000,
31'b1000100000000010000000000000000,
31'b0000000000000100000000000000000,
31'b0000000001000100000000000000000,
31'b0010000000000001000000000000000,
31'b1001000000000000000000000001000,
31'b0000000100000100000000000000000,
31'b0000001000000000000001000000000,
31'b0000100000000000000000100000010,
31'b0100000000100000000000000100000,
31'b0000001000000100000000000000000,
31'b0000000100000000000001000000000,
31'b0000010000000000001000000000000,
31'b0000000010000000000001000000000,
31'b0000000001000000000001000000000,
31'b0000000000000000000001000000000,
31'b0100000000010000000000000010000,
31'b1100000000000000010000000000000,
31'b0000010000000100000000000000000,
31'b0110000000000000000000100000000,
31'b0000001000000000001000000000000,
31'b0001000000000001010000000000000,
31'b0000000000000000000000100001000,
31'b0000011000000000000001000000000,
31'b0000000100000000001000000000000,
31'b1000000000000001000000010000000,
31'b1000000000010000000000000000000,
31'b0000000000000000010000000010000,
31'b0000000000000000001000000000000,
31'b0000000001000000001000000000000,
31'b0000000010000000001000000000000,
31'b0000010000000000000001000000000,
31'b0000000000000000000000010100000,
31'b1000000000000010000000000000000,
31'b0000100000000100000000000000000,
31'b1000000010000010000000000000000,
31'b0100000000000000000100000010000,
31'b1000000100000010000000000000000,
31'b1000001000000000000100000000000,
31'b0000000000001000000000000010000,
31'b0000000000000000000000100000010,
31'b0010000000000000000000000000001,
31'b1000000100000000000100000000000,
31'b1000000000000000000000010000100,
31'b1000000010000000000100000000000,
31'b1100000000001000000000000000000,
31'b1000000000000000000100000000000,
31'b0000100000000000000001000000000,
31'b1000000000000000000000001010000,
31'b0000000000000000100000100000000,
31'b0100001000000000000000001000000,
31'b0100000000000000000000000001100,
31'b0001000000100000000000000000000,
31'b0001000001100000000000000000000,
31'b0010000000000000000000000000100,
31'b1100000000000000000010000000000,
31'b0100000010000000000000001000000,
31'b0010010000000000000000000000001,
31'b0100000000000000000000001000000,
31'b1001000000000000000000000000010,
31'b0000100000000000001000000000000,
31'b0000000000000000000010000010000,
31'b1000010000000000000100000000000,
31'b0100000000000001000000000000010
};

parameter [0:31*(2**15)-1] SYNDROME_TABLE_31_16 = {
31'b0000000000000000000000000000000,
31'b0000000000000010000000000000000,
31'b0000000000000100000000000000000,
31'b0000000000000110000000000000000,
31'b0000000000001000000000000000000,
31'b0000000000001010000000000000000,
31'b0000000000001100000000000000000,
31'b0000000000001110000000000000000,
31'b0000000000010000000000000000000,
31'b0000000000010010000000000000000,
31'b0000000000010100000000000000000,
31'b0000000000010110000000000000000,
31'b0000000000011000000000000000000,
31'b0000000000011010000000000000000,
31'b0000000000011100000000000000000,
31'b0011001000000000001000000000000,
31'b0000000000100000000000000000000,
31'b0000000000100010000000000000000,
31'b0000000000100100000000000000000,
31'b0000000000100110000000000000000,
31'b0000000000101000000000000000000,
31'b0000000000101010000000000000000,
31'b0000000000101100000000000000000,
31'b0001000000000000010000010000100,
31'b0000000000110000000000000000000,
31'b0000000000110010000000000000000,
31'b0000000000110100000000000000000,
31'b0000010000000000001010000000100,
31'b0000000000111000000000000000000,
31'b0100001000000000000010010000000,
31'b0110010000000000010000000000000,
31'b0110010000000010010000000000000,
31'b0000000001000000000000000000000,
31'b0000000001000010000000000000000,
31'b0000000001000100000000000000000,
31'b0000000001000110000000000000000,
31'b0000000001001000000000000000000,
31'b0000000001001010000000000000000,
31'b0000000001001100000000000000000,
31'b0001000000000000000000000011000,
31'b0000000001010000000000000000000,
31'b0000000001010010000000000000000,
31'b0000000001010100000000000000000,
31'b0000000001010110000000000000000,
31'b0000000001011000000000000000000,
31'b0000001000000000100000000100000,
31'b0010000000000000100000100001000,
31'b0001000000010000000000000011000,
31'b0000000001100000000000000000000,
31'b0000000001100010000000000000000,
31'b0000000001100100000000000000000,
31'b0000000100000000000100000010100,
31'b0000000001101000000000000000000,
31'b0000100100000000000000010000000,
31'b0000100000000000010100000001000,
31'b0001000000100000000000000011000,
31'b0000000001110000000000000000000,
31'b1000000100000000000010000100000,
31'b1000010000000000000100100000000,
31'b1000010000000010000100100000000,
31'b1100100000000000100000000000000,
31'b0000100100010000000000010000000,
31'b1100100000000100100000000000000,
31'b0001001000000000000001010000010,
31'b0000000010000000000000000000000,
31'b0000000010000010000000000000000,
31'b0000000010000100000000000000000,
31'b0000000010000110000000000000000,
31'b0000000010001000000000000000000,
31'b0000000010001010000000000000000,
31'b0000000010001100000000000000000,
31'b0001000000000000100000100100000,
31'b0000000010010000000000000000000,
31'b0000000010010010000000000000000,
31'b0000000010010100000000000000000,
31'b0000000000000000101000000001000,
31'b0000000010011000000000000000000,
31'b0000001000000000000000100011000,
31'b0010000000000000000000000110000,
31'b0010000000000010000000000110000,
31'b0000000010100000000000000000000,
31'b0000000010100010000000000000000,
31'b0000000010100100000000000000000,
31'b0000000010100110000000000000000,
31'b0000000010101000000000000000000,
31'b0000000010101010000000000000000,
31'b0000000010101100000000000000000,
31'b0001000010000000010000010000100,
31'b0000000010110000000000000000000,
31'b0000000010110010000000000000000,
31'b0000010000000001000000001000000,
31'b0000010000000011000000001000000,
31'b0100000000000001000001000010000,
31'b0100001010000000000010010000000,
31'b0010000000100000000000000110000,
31'b1010010000000000001100000000000,
31'b0000000011000000000000000000000,
31'b0000000011000010000000000000000,
31'b0000000011000100000000000000000,
31'b0010001000000000100000000010000,
31'b0000000011001000000000000000000,
31'b0010000000000000001000100000000,
31'b0000001000000000001000000101000,
31'b0010000000000100001000100000000,
31'b0000000011010000000000000000000,
31'b0011000000000000000000000101000,
31'b0001001000000000000000100000000,
31'b0001001000000010000000100000000,
31'b0001000000000000101000000010000,
31'b0010000000010000001000100000000,
31'b0010000001000000000000000110000,
31'b0010000001000010000000000110000,
31'b0000000011100000000000000000000,
31'b0010000100000000000000000000011,
31'b0000001000000000000100001000001,
31'b0010001000100000100000000010000,
31'b0000100000000000001001000000001,
31'b0010000000100000001000100000000,
31'b0000100010000000010100000001000,
31'b1100100000000000001000000001000,
31'b1001000000000001000000000000001,
31'b1001000000000011000000000000001,
31'b0001001000100000000000100000000,
31'b0101000000000001000001000001000,
31'b1100100010000000100000000000000,
31'b0010000100000000000100000100100,
31'b0010010000000000000010100000100,
31'b1100010000000001000010000000000,
31'b0000000100000000000000000000000,
31'b0000000100000010000000000000000,
31'b0000000100000100000000000000000,
31'b0000000100000110000000000000000,
31'b0000000100001000000000000000000,
31'b0000000100001010000000000000000,
31'b0000000100001100000000000000000,
31'b0001100000000001000100000000000,
31'b0000000100010000000000000000000,
31'b0000000100010010000000000000000,
31'b0000000100010100000000000000000,
31'b1000000000000000001101000000000,
31'b0000000100011000000000000000000,
31'b1000101000000000000000001000000,
31'b0010000000000001000001001000000,
31'b1000101000000100000000001000000,
31'b0000000100100000000000000000000,
31'b0000000100100010000000000000000,
31'b0000000100100100000000000000000,
31'b0000000100100110000000000000000,
31'b0000000100101000000000000000000,
31'b0000100001000000000000010000000,
31'b0000000000000001010000000010000,
31'b0000100001000100000000010000000,
31'b0000000100110000000000000000000,
31'b1000000001000000000010000100000,
31'b0000010000000000000001000110000,
31'b1000000001000100000010000100000,
31'b0100000000000000000000001100000,
31'b0100000000000010000000001100000,
31'b0100000000000100000000001100000,
31'b0100000000000110000000001100000,
31'b0000000101000000000000000000000,
31'b0000000101000010000000000000000,
31'b0000000101000100000000000000000,
31'b0000000101000110000000000000000,
31'b0000000101001000000000000000000,
31'b0000100000100000000000010000000,
31'b0000000101001100000000000000000,
31'b0001000100000000000000000011000,
31'b0000000101010000000000000000000,
31'b1000000000100000000010000100000,
31'b0000000101010100000000000000000,
31'b1000000001000000001101000000000,
31'b0000000101011000000000000000000,
31'b0000100000110000000000010000000,
31'b0010000100000000100000100001000,
31'b0001111000000000000000000000001,
31'b0000000101100000000000000000000,
31'b0000100000001000000000010000000,
31'b0000000101100100000000000000000,
31'b0000000000000000000100000010100,
31'b0000100000000010000000010000000,
31'b0000100000000000000000010000000,
31'b0000100000000110000000010000000,
31'b0000100000000100000000010000000,
31'b1000000000000010000010000100000,
31'b1000000000000000000010000100000,
31'b1000010100000000000100100000000,
31'b1000000000000100000010000100000,
31'b0100000001000000000000001100000,
31'b0000100000010000000000010000000,
31'b0100100000000000011000000000001,
31'b0000100000010100000000010000000,
31'b0000000110000000000000000000000,
31'b0000000110000010000000000000000,
31'b0000000110000100000000000000000,
31'b0100000000000000100100000000001,
31'b0000000110001000000000000000000,
31'b0000110000000000000000100000001,
31'b0100010000000001000000000100000,
31'b0100010000000011000000000100000,
31'b0000000110010000000000000000000,
31'b1000000000000000010000000001001,
31'b0100000000000000010001000000000,
31'b0100000000000010010001000000000,
31'b0000010000000000010000001010000,
31'b1000101010000000000000001000000,
31'b0100000000001000010001000000000,
31'b0100000000001010010001000000000,
31'b0000000110100000000000000000000,
31'b0010000001000000000000000000011,
31'b0110000000000000000000001010000,
31'b0110000000000010000000001010000,
31'b0010010000000000000001000000000,
31'b0010010000000010000001000000000,
31'b0010010000000100000001000000000,
31'b1010000001000000000010000010000,
31'b0010000000000001010000000100000,
31'b1000000011000000000010000100000,
31'b0100000000100000010001000000000,
31'b0101000000000000100000101000000,
31'b0100000010000000000000001100000,
31'b0101000000000000000001010000100,
31'b0100000010000100000000001100000,
31'b1000100001000000000100000000001,
31'b0000000111000000000000000000000,
31'b0010000000100000000000000000011,
31'b0100001000000000000000000000110,
31'b0100001000000010000000000000110,
31'b0000010000000000001000010000010,
31'b0010000100000000001000100000000,
31'b0100010001000001000000000100000,
31'b1010000000100000000010000010000,
31'b0001000000000000010010000000010,
31'b1000000010100000000010000100000,
31'b0100000001000000010001000000000,
31'b0100011000000001100000000000000,
31'b0001000100000000101000000010000,
31'b0010000100010000001000100000000,
31'b1010000000000000000101100000000,
31'b1000100000100000000100000000001,
31'b0010000000000010000000000000011,
31'b0010000000000000000000000000011,
31'b0110000001000000000000001010000,
31'b0010000000000100000000000000011,
31'b0010010001000000000001000000000,
31'b0000100010000000000000010000000,
31'b1010000000000010000010000010000,
31'b1010000000000000000010000010000,
31'b1001000100000001000000000000001,
31'b1000000010000000000010000100000,
31'b0100001000000000001000001001000,
31'b1000100000001000000100000000001,
31'b0100100000000000000101000001000,
31'b0010000000000000000100000100100,
31'b1001000000000000100010100000000,
31'b1000100000000000000100000000001,
31'b0000001000000000000000000000000,
31'b0000001000000010000000000000000,
31'b0000001000000100000000000000000,
31'b0000001000000110000000000000000,
31'b0000001000001000000000000000000,
31'b0000001000001010000000000000000,
31'b0000001000001100000000000000000,
31'b0011000000010000001000000000000,
31'b0000001000010000000000000000000,
31'b0000001000010010000000000000000,
31'b0000001000010100000000000000000,
31'b0011000000001000001000000000000,
31'b0000001000011000000000000000000,
31'b0000000001000000100000000100000,
31'b0011000000000010001000000000000,
31'b0011000000000000001000000000000,
31'b0000001000100000000000000000000,
31'b0000001000100010000000000000000,
31'b0000001000100100000000000000000,
31'b0110000000000000000000000000101,
31'b0000001000101000000000000000000,
31'b0100000000010000000010010000000,
31'b0000001000101100000000000000000,
31'b0110000000001000000000000000101,
31'b0000001000110000000000000000000,
31'b0100000000001000000010010000000,
31'b0001010000000000000000010000001,
31'b0110000000010000000000000000101,
31'b0100000000000010000010010000000,
31'b0100000000000000000010010000000,
31'b0110011000000000010000000000000,
31'b0100000000000100000010010000000,
31'b0000001001000000000000000000000,
31'b0000001001000010000000000000000,
31'b0000001001000100000000000000000,
31'b0010000010000000100000000010000,
31'b0000001001001000000000000000000,
31'b0000000000010000100000000100000,
31'b0000001001001100000000000000000,
31'b0001001000000000000000000011000,
31'b0000001001010000000000000000000,
31'b0000000000001000100000000100000,
31'b0001000010000000000000100000000,
31'b0001000010000010000000100000000,
31'b0000000000000010100000000100000,
31'b0000000000000000100000000100000,
31'b0001000010001000000000100000000,
31'b0000000000000100100000000100000,
31'b0000001001100000000000000000000,
31'b0100000100000000100000001000000,
31'b0000001001100100000000000000000,
31'b0110000001000000000000000000101,
31'b0000100000000000000010001100000,
31'b0000101100000000000000010000000,
31'b0000101000000000010100000001000,
31'b0001001000100000000000000011000,
31'b1000000000000000000000011000000,
31'b1000000000000010000000011000000,
31'b1000000000000100000000011000000,
31'b1000000000000110000000011000000,
31'b1000000000001000000000011000000,
31'b0000000000100000100000000100000,
31'b1000000000001100000000011000000,
31'b0001000000000000000001010000010,
31'b0000001010000000000000000000000,
31'b0000001010000010000000000000000,
31'b0000001010000100000000000000000,
31'b0010000001000000100000000010000,
31'b0000001010001000000000000000000,
31'b0000001010001010000000000000000,
31'b0000001010001100000000000000000,
31'b0011000010010000001000000000000,
31'b0000001010010000000000000000000,
31'b0000001010010010000000000000000,
31'b0001000001000000000000100000000,
31'b0001000001000010000000100000000,
31'b0000001010011000000000000000000,
31'b0000000000000000000000100011000,
31'b0010001000000000000000000110000,
31'b0011000010000000001000000000000,
31'b0000001010100000000000000000000,
31'b0100000000000000000100000010010,
31'b0000001010100100000000000000000,
31'b0110000010000000000000000000101,
31'b0000001010101000000000000000000,
31'b0100000010010000000010010000000,
31'b0000001010101100000000000000000,
31'b1100000000000000000110000000001,
31'b0000001010110000000000000000000,
31'b0100000010001000000010010000000,
31'b0001000001100000000000100000000,
31'b0001010100000000001001000000000,
31'b0100001000000001000001000010000,
31'b0100000010000000000010010000000,
31'b0011110000000000000000000000010,
31'b1110100000000000000000000010000,
31'b0000001011000000000000000000000,
31'b0010000000000100100000000010000,
31'b0001000000010000000000100000000,
31'b0010000000000000100000000010000,
31'b0000001011001000000000000000000,
31'b0010001000000000001000100000000,
31'b0000000000000000001000000101000,
31'b0010000000001000100000000010000,
31'b0001000000000100000000100000000,
31'b0001000000000110000000100000000,
31'b0001000000000000000000100000000,
31'b0001000000000010000000100000000,
31'b0001000000001100000000100000000,
31'b0000000010000000100000000100000,
31'b0001000000001000000000100000000,
31'b0001000000001010000000100000000,
31'b0000001011100000000000000000000,
31'b0100000110000000100000001000000,
31'b0000000000000000000100001000001,
31'b0010000000100000100000000010000,
31'b0000101000000000001001000000001,
31'b0010001000100000001000100000000,
31'b0000000000100000001000000101000,
31'b1010000000000001001000000000001,
31'b1000000010000000000000011000000,
31'b1001000000000000000001000100100,
31'b0001000000100000000000100000000,
31'b0001000000100010000000100000000,
31'b1001000000000000110000000000010,
31'b0000000010100000100000000100000,
31'b0001000000101000000000100000000,
31'b0001000010000000000001010000010,
31'b0000001100000000000000000000000,
31'b0000001100000010000000000000000,
31'b0000001100000100000000000000000,
31'b0010000000000000000100001000010,
31'b0000001100001000000000000000000,
31'b1000100000010000000000001000000,
31'b1000000000000001001000000000010,
31'b1000100000010100000000001000000,
31'b0000001100010000000000000000000,
31'b1000100000001000000000001000000,
31'b0001100000000000000001000000010,
31'b1000100000001100000000001000000,
31'b1000100000000010000000001000000,
31'b1000100000000000000000001000000,
31'b1000100000000110000000001000000,
31'b1000100000000100000000001000000,
31'b0000001100100000000000000000000,
31'b0100000001000000100000001000000,
31'b0000001100100100000000000000000,
31'b0110000100000000000000000000101,
31'b1000000000000000100010000000000,
31'b1000000000000010100010000000000,
31'b1000000000000100100010000000000,
31'b1000110010000001000000000000000,
31'b0000100000000000100000010100000,
31'b1000100000101000000000001000000,
31'b0001100000100000000001000000010,
31'b0011000000000000000000100000011,
31'b1000000000010000100010000000000,
31'b1000100000100000000000001000000,
31'b1000000000010100100010000000000,
31'b1000100000100100000000001000000,
31'b0000001101000000000000000000000,
31'b0100000000100000100000001000000,
31'b0100000010000000000000000000110,
31'b0100000010000010000000000000110,
31'b1100000000000000000000010100000,
31'b0000101000100000000000010000000,
31'b1100000000000100000000010100000,
31'b0001110000010000000000000000001,
31'b0100100000000000000010000000000,
31'b0100100000000010000010000000000,
31'b0100100000000100000010000000000,
31'b0100100000000110000010000000000,
31'b0100100000001000000010000000000,
31'b0000000100000000100000000100000,
31'b0100100000001100000010000000000,
31'b0001110000000000000000000000001,
31'b0100000000000010100000001000000,
31'b0100000000000000100000001000000,
31'b0100000010100000000000000000110,
31'b0100000000000100100000001000000,
31'b1000000001000000100010000000000,
31'b0000101000000000000000010000000,
31'b1010000000000001000001010000000,
31'b0000101000000100000000010000000,
31'b1000000100000000000000011000000,
31'b1000001000000000000010000100000,
31'b1010000000000000000010100001000,
31'b1000001000000100000010000100000,
31'b1000000100001000000000011000000,
31'b0000101000010000000000010000000,
31'b0011010000000000000001100000000,
31'b0001110000100000000000000000001,
31'b0000001110000000000000000000000,
31'b0000001110000010000000000000000,
31'b0100000001000000000000000000110,
31'b0100001000000000100100000000001,
31'b1000010000000000000000000001100,
31'b1000100010010000000000001000000,
31'b1000010000000100000000000001100,
31'b1000110000100001000000000000000,
31'b0000100000000000010000100000100,
31'b1000100010001000000000001000000,
31'b0100001000000000010001000000000,
31'b0100010001000001100000000000000,
31'b1000100010000010000000001000000,
31'b1000100010000000000000001000000,
31'b0100001000001000010001000000000,
31'b1000100010000100000000001000000,
31'b0010000000000000100100000000100,
31'b0100000100000000000100000010010,
31'b0110001000000000000000001010000,
31'b1001000000000000000010100100000,
31'b1000000010000000100010000000000,
31'b1000110000000101000000000000000,
31'b1000110000000011000000000000000,
31'b1000110000000001000000000000000,
31'b0010001000000001010000000100000,
31'b0010010000000001000100000000010,
31'b0100001000100000010001000000000,
31'b0001010000000000001001000000000,
31'b1000010000000000001000001000010,
31'b1000100010100000000000001000000,
31'b1000100000000000100000000000110,
31'b1000000000000000001010000001000,
31'b0100000000000100000000000000110,
31'b0100000010100000100000001000000,
31'b0100000000000000000000000000110,
31'b0100000000000010000000000000110,
31'b1100000010000000000000010100000,
31'b0010001100000000001000100000000,
31'b0100000000001000000000000000110,
31'b0100000000001010000000000000110,
31'b0100100010000000000010000000000,
31'b0100100010000010000010000000000,
31'b0001000100000000000000100000000,
31'b0100010000000001100000000000000,
31'b0100100010001000000010000000000,
31'b0000100000000001000100100000000,
31'b0100000000000000000100000100001,
31'b0100010000001001100000000000000,
31'b0100000010000010100000001000000,
31'b0100000010000000100000001000000,
31'b0100000000100000000000000000110,
31'b0100000010000100100000001000000,
31'b1000010000000000010000010010000,
31'b0010000000000001110000000000000,
31'b0101000000000000000000101100000,
31'b1010001000000000000010000010000,
31'b1001000000000000001010000010000,
31'b1000001010000000000010000100000,
31'b0100000000000000001000001001000,
31'b0100010000100001100000000000000,
31'b0010010000000000010000000000110,
31'b0010001000000000000100000100100,
31'b0001000000000000001000000000011,
31'b1000101000000000000100000000001,
31'b0000010000000000000000000000000,
31'b0000010000000010000000000000000,
31'b0000010000000100000000000000000,
31'b0000010000000110000000000000000,
31'b0000010000001000000000000000000,
31'b0000010000001010000000000000000,
31'b0000010000001100000000000000000,
31'b0101000000000000000010000000001,
31'b0000010000010000000000000000000,
31'b0000010000010010000000000000000,
31'b0000010000010100000000000000000,
31'b0000010000010110000000000000000,
31'b0000010000011000000000000000000,
31'b0000010000011010000000000000000,
31'b0110000000100000010000000000000,
31'b0110000000100010010000000000000,
31'b0000010000100000000000000000000,
31'b0000010000100010000000000000000,
31'b0000010000100100000000000000000,
31'b0000010000100110000000000000000,
31'b0000010000101000000000000000000,
31'b0010000000000000001000010000001,
31'b0110000000010000010000000000000,
31'b0110000000010010010000000000000,
31'b0000010000110000000000000000000,
31'b0000010000110010000000000000000,
31'b0000000010000001000000001000000,
31'b0000000000000000001010000000100,
31'b0110000000000100010000000000000,
31'b0110000000000110010000000000000,
31'b0110000000000000010000000000000,
31'b0110000000000010010000000000000,
31'b0000010001000000000000000000000,
31'b0000010001000010000000000000000,
31'b0000010001000100000000000000000,
31'b1000000000000000000011000010000,
31'b0000010001001000000000000000000,
31'b0000000000000000000001000000011,
31'b1100000000000000000000000001010,
31'b0001010000000000000000000011000,
31'b0000010001010000000000000000000,
31'b0000010001010010000000000000000,
31'b1000000000100000000100100000000,
31'b1000000000100010000100100000000,
31'b0000010001011000000000000000000,
31'b0000011000000000100000000100000,
31'b1100000000010000000000000001010,
31'b0001101100000000000000000000001,
31'b0000010001100000000000000000000,
31'b0000010001100010000000000000000,
31'b1000000000010000000100100000000,
31'b1000000000100000000011000010000,
31'b0010100000000000000000100000010,
31'b0000110100000000000000010000000,
31'b1100000000100000000000000001010,
31'b0001010000100000000000000011000,
31'b1000000000000100000100100000000,
31'b1000010100000000000010000100000,
31'b1000000000000000000100100000000,
31'b1000000000000010000100100000000,
31'b1100110000000000100000000000000,
31'b0001100000000000100000000010010,
31'b1000000000001000000100100000000,
31'b1100000010000001000010000000000,
31'b0000010010000000000000000000000,
31'b0000010010000010000000000000000,
31'b0000010010000100000000000000000,
31'b0000100000000001100010000000000,
31'b0000010010001000000000000000000,
31'b0000100100000000000000100000001,
31'b0100000100000001000000000100000,
31'b0101000010000000000010000000001,
31'b0000010010010000000000000000000,
31'b0000100000000000000000001001100,
31'b0000000000100001000000001000000,
31'b0000010000000000101000000001000,
31'b0000010010011000000000000000000,
31'b0000100100010000000000100000001,
31'b0010010000000000000000000110000,
31'b1010000000100000001100000000000,
31'b0000010010100000000000000000000,
31'b0000100000000000001000000000010,
31'b0000000000010001000000001000000,
31'b0000100000000100001000000000010,
31'b0010000100000000000001000000000,
31'b0010000100000010000001000000000,
31'b0010000100000100000001000000000,
31'b1010000000010000001100000000000,
31'b0000000000000101000000001000000,
31'b0000100000010000001000000000010,
31'b0000000000000001000000001000000,
31'b0000000000000011000000001000000,
31'b0010000100010000000001000000000,
31'b1010000000000100001100000000000,
31'b0000000000001001000000001000000,
31'b1010000000000000001100000000000,
31'b0000010011000000000000000000000,
31'b0010100000000000000001010000000,
31'b1000001000000001000000010000000,
31'b1000001000000011000000010000000,
31'b0000010011001000000000000000000,
31'b0010010000000000001000100000000,
31'b1100000010000000000000000001010,
31'b0010010000000100001000100000000,
31'b0001000000000000000100011000000,
31'b0011010000000000000000000101000,
31'b0001011000000000000000100000000,
31'b0100001100000001100000000000000,
31'b0001010000000000101000000010000,
31'b1100000000000000101000000000010,
31'b0010010001000000000000000110000,
31'b1100000000100001000010000000000,
31'b0000000000000000000000110000001,
31'b0000100001000000001000000000010,
31'b0000000001010001000000001000000,
31'b0100100000000001000000010100000,
31'b0010000101000000000001000000000,
31'b0010010000100000001000100000000,
31'b0010000101000100000001000000000,
31'b1100000000010001000010000000000,
31'b0000000001000101000000001000000,
31'b0100000000000100011000100000000,
31'b0000000001000001000000001000000,
31'b0100000000000000011000100000000,
31'b0010000101010000000001000000000,
31'b1100000000000101000010000000000,
31'b0010000000000000000010100000100,
31'b1100000000000001000010000000000,
31'b0000010100000000000000000000000,
31'b0000010100000010000000000000000,
31'b0000010100000100000000000000000,
31'b0000010100000110000000000000000,
31'b0000010100001000000000000000000,
31'b0000100010000000000000100000001,
31'b0100000010000001000000000100000,
31'b0101000100000000000010000000001,
31'b0000010100010000000000000000000,
31'b1000000000000000000000100010100,
31'b0000010100010100000000000000000,
31'b1000010000000000001101000000000,
31'b0000010100011000000000000000000,
31'b1000111000000000000000001000000,
31'b0110000100100000010000000000000,
31'b1000100000000000000100110000000,
31'b0000010100100000000000000000000,
31'b0000010100100010000000000000000,
31'b0000010100100100000000000000000,
31'b0000010100100110000000000000000,
31'b0010000010000000000001000000000,
31'b0010000010000010000001000000000,
31'b0010000010000100000001000000000,
31'b1010000000000000110000010000000,
31'b0000010100110000000000000000000,
31'b1000010001000000000010000100000,
31'b0000000000000000000001000110000,
31'b0000000100000000001010000000100,
31'b0100010000000000000000001100000,
31'b0110000000000000000100010001000,
31'b0110000100000000010000000000000,
31'b0110000100000010010000000000000,
31'b0000010101000000000000000000000,
31'b0000010101000010000000000000000,
31'b1000000000000000001000000100100,
31'b1000000100000000000011000010000,
31'b0000010101001000000000000000000,
31'b0000110000100000000000010000000,
31'b1100000100000000000000000001010,
31'b0001101000010000000000000000001,
31'b0000010101010000000000000000000,
31'b1000010000100000000010000100000,
31'b1000000100100000000100100000000,
31'b0110100000000000010000010000000,
31'b0000010101011000000000000000000,
31'b0001101000000100000000000000001,
31'b1001000000000000000000100001100,
31'b0001101000000000000000000000001,
31'b0000010101100000000000000000000,
31'b0000000000000000001001100000000,
31'b1000000100010000000100100000000,
31'b0000010000000000000100000010100,
31'b0010000011000000000001000000000,
31'b0000110000000000000000010000000,
31'b0010101000000000010010000000000,
31'b0000110000000100000000010000000,
31'b1000010000000010000010000100000,
31'b1000010000000000000010000100000,
31'b1000000100000000000100100000000,
31'b1000010000000100000010000100000,
31'b0111100000000000000000000000100,
31'b0001000000000000000001000101000,
31'b1101000000000000000000000100001,
31'b0001101000100000000000000000001,
31'b0000010110000000000000000000000,
31'b0000100000001000000000100000001,
31'b0100000000001001000000000100000,
31'b0100010000000000100100000000001,
31'b0010000000100000000001000000000,
31'b0000100000000000000000100000001,
31'b0100000000000001000000000100000,
31'b0100000000000011000000000100000,
31'b0000010110010000000000000000000,
31'b1000010000000000010000000001001,
31'b0100010000000000010001000000000,
31'b0100010000000010010001000000000,
31'b0000000000000000010000001010000,
31'b0000100000010000000000100000001,
31'b0100000000010001000000000100000,
31'b0100000001000000010000000000011,
31'b0010000000001000000001000000000,
31'b0010000000001010000001000000000,
31'b0010000000001100000001000000000,
31'b1011000000000000000000001000010,
31'b0010000000000000000001000000000,
31'b0010000000000010000001000000000,
31'b0010000000000100000001000000000,
31'b1000101000000001000000000000000,
31'b0010000000011000000001000000000,
31'b0010001000000001000100000000010,
31'b0000000100000001000000001000000,
31'b0001001000000000001001000000000,
31'b0010000000010000000001000000000,
31'b0010000000010010000001000000000,
31'b0010000000010100000001000000000,
31'b1010000100000000001100000000000,
31'b0000010111000000000000000000000,
31'b0010100100000000000001010000000,
31'b1000001100000001000000010000000,
31'b1001001000000000000000000010100,
31'b0000000000000000001000010000010,
31'b0000100001000000000000100000001,
31'b0100000001000001000000000100000,
31'b0100000001000011000000000100000,
31'b0001010000000000010010000000010,
31'b1100000000000000010010000010000,
31'b0100010001000000010001000000000,
31'b0100001000000001100000000000000,
31'b0000000001000000010000001010000,
31'b0100000000000100010000000000011,
31'b0100000001010001000000000100000,
31'b0100000000000000010000000000011,
31'b0010000001001000000001000000000,
31'b0010010000000000000000000000011,
31'b0010000001001100000001000000000,
31'b0011000000000000000001000011000,
31'b0010000001000000000001000000000,
31'b0010000001000010000001000000000,
31'b0010000001000100000001000000000,
31'b1010010000000000000010000010000,
31'b0010000001011000000001000000000,
31'b1100000000000000100000100000001,
31'b0000000101000001000000001000000,
31'b0100001000100001100000000000000,
31'b0010000001010000000001000000000,
31'b0010010000000000000100000100100,
31'b0010000100000000000010100000100,
31'b1100000100000001000010000000000,
31'b0000011000000000000000000000000,
31'b0000011000000010000000000000000,
31'b0000011000000100000000000000000,
31'b0010000000000000010010010000000,
31'b0000011000001000000000000000000,
31'b0000011000001010000000000000000,
31'b0100000000000000001000010000100,
31'b0101001000000000000010000000001,
31'b0000011000010000000000000000000,
31'b0000011000010010000000000000000,
31'b0001000000100000000000010000001,
31'b0011010000001000001000000000000,
31'b0000011000011000000000000000000,
31'b0000000000000000010000000000101,
31'b0110001000100000010000000000000,
31'b0011010000000000001000000000000,
31'b0000011000100000000000000000000,
31'b0101000000000000011000000000000,
31'b0001000000010000000000010000001,
31'b0110010000000000000000000000101,
31'b0011000000000000000010000000100,
31'b0101000000001000011000000000000,
31'b0110001000010000010000000000000,
31'b1000100110000001000000000000000,
31'b0001000000000100000000010000001,
31'b0101000000010000011000000000000,
31'b0001000000000000000000010000001,
31'b0001000000000010000000010000001,
31'b0110001000000100010000000000000,
31'b0100010000000000000010010000000,
31'b0110001000000000010000000000000,
31'b0110001000000010010000000000000,
31'b0000011001000000000000000000000,
31'b0000011001000010000000000000000,
31'b1000000010000001000000010000000,
31'b1000001000000000000011000010000,
31'b0000011001001000000000000000000,
31'b0000010000010000100000000100000,
31'b1100001000000000000000000001010,
31'b0001100100010000000000000000001,
31'b0000000000000001000100000000001,
31'b0000010000001000100000000100000,
31'b0001010010000000000000100000000,
31'b0100100000000000000100100100000,
31'b0000010000000010100000000100000,
31'b0000010000000000100000000100000,
31'b0001100100000010000000000000001,
31'b0001100100000000000000000000001,
31'b0001000000000001000000101000000,
31'b0101000001000000011000000000000,
31'b1000001000010000000100100000000,
31'b0110000000000000110000000100000,
31'b0011000001000000000010000000100,
31'b0000111100000000000000010000000,
31'b0110000000000000000001000000110,
31'b0000100000000000000000000101010,
31'b1000010000000000000000011000000,
31'b1010000000000000000100000101000,
31'b1000001000000000000100100000000,
31'b1000001000000010000100100000000,
31'b1000010000001000000000011000000,
31'b0000010000100000100000000100000,
31'b1100000000000000000001010010000,
31'b0001100100100000000000000000001,
31'b0000011010000000000000000000000,
31'b1000100000000000010000000010000,
31'b1000000001000001000000010000000,
31'b1000100000000100010000000010000,
31'b1000000100000000000000000001100,
31'b1000100000001000010000000010000,
31'b1000000100000100000000000001100,
31'b1000100100100001000000000000000,
31'b1000000000000000000000101000001,
31'b1000100000010000010000000010000,
31'b0001010001000000000000100000000,
31'b0100000101000001100000000000000,
31'b1000000100010000000000000001100,
31'b0000010000000000000000100011000,
31'b0011100000100000000000000000010,
31'b0011010010000000001000000000000,
31'b1001000000000000000100000000000,
31'b1001000000000010000100000000000,
31'b1001000000000100000100000000000,
31'b1001000000000110000100000000000,
31'b1001000000001000000100000000000,
31'b1001000000001010000100000000000,
31'b1001000000001100000100000000000,
31'b1000100100000001000000000000000,
31'b1001000000010000000100000000000,
31'b1010100000000000000001001000000,
31'b0000001000000001000000001000000,
31'b0001000100000000001001000000000,
31'b1001000000011000000100000000000,
31'b0100010010000000000010010000000,
31'b0011100000000000000000000000010,
31'b1010001000000000001100000000000,
31'b1000000000000101000000010000000,
31'b1000100001000000010000000010000,
31'b1000000000000001000000010000000,
31'b1000000000000011000000010000000,
31'b1000000101000000000000000001100,
31'b0110000000000000100001001000000,
31'b1000000000001001000000010000000,
31'b1000000000100000000100000011000,
31'b0001010000000100000000100000000,
31'b0100000100000101100000000000000,
31'b0001010000000000000000100000000,
31'b0100000100000001100000000000000,
31'b0101100000000000100100000000000,
31'b0100000000000000000010100000001,
31'b0001010000001000000000100000000,
31'b0100000100001001100000000000000,
31'b1001000001000000000100000000000,
31'b1001000001000010000100000000000,
31'b1000000000100001000000010000000,
31'b1000000000100011000000010000000,
31'b1001000001001000000100000000000,
31'b1001000000000001010000000000100,
31'b1000000000101001000000010000000,
31'b1000000000000000000100000011000,
31'b1001000001010000000100000000000,
31'b0100000100000000001010000000010,
31'b0001010000100000000000100000000,
31'b0100001000000000011000100000000,
31'b0110100000000000000011000000000,
31'b0100000000000000110000000010000,
31'b0011100001000000000000000000010,
31'b1100001000000001000010000000000,
31'b0000011100000000000000000000000,
31'b0000011100000010000000000000000,
31'b0000011100000100000000000000000,
31'b0010010000000000000100001000010,
31'b1000000010000000000000000001100,
31'b1000110000010000000000001000000,
31'b1000010000000001001000000000010,
31'b1000100010100001000000000000000,
31'b0000100000000000000000000011001,
31'b1000110000001000000000001000000,
31'b0001110000000000000001000000010,
31'b1100100000000000000001000010000,
31'b1000110000000010000000001000000,
31'b1000110000000000000000001000000,
31'b1000100000000000000010000001010,
31'b1000000000000000101000000000100,
31'b0001000000000000100001000001000,
31'b0101000100000000011000000000000,
31'b0001000100010000000000010000001,
31'b1101000000000000100000000000001,
31'b1000010000000000100010000000000,
31'b1000100010000101000000000000000,
31'b1000100010000011000000000000000,
31'b1000100010000001000000000000000,
31'b0001000100000100000000010000001,
31'b0010000010000001000100000000010,
31'b0001000100000000000000010000001,
31'b0001000010000000001001000000000,
31'b1000010000010000100010000000000,
31'b1000110000100000000000001000000,
31'b0110001100000000010000000000000,
31'b1000100010010001000000000000000,
31'b0100000000000001001000000001000,
31'b0100010000100000100000001000000,
31'b1000001000000000001000000100100,
31'b1001000010000000000000000010100,
31'b1100010000000000000000010100000,
31'b0001100000010100000000000000001,
31'b0010100000100000010010000000000,
31'b0001100000010000000000000000001,
31'b0100110000000000000010000000000,
31'b0100110000000010000010000000000,
31'b0100110000000100000010000000000,
31'b0100000010000001100000000000000,
31'b0101000000000001000000100100000,
31'b0001100000000100000000000000001,
31'b0001100000000010000000000000001,
31'b0001100000000000000000000000001,
31'b0100010000000010100000001000000,
31'b0100010000000000100000001000000,
31'b0100100000000010001000000000100,
31'b0100100000000000001000000000100,
31'b1000010001000000100010000000000,
31'b0000111000000000000000010000000,
31'b0010100000000000010010000000000,
31'b0000000000000000100001000010000,
31'b1000010100000000000000011000000,
31'b1010000000000000000000101000010,
31'b1010000000000000010000010100000,
31'b0100100000010000001000000000100,
31'b0011000000000100000001100000000,
31'b0001100000100100000000000000001,
31'b0011000000000000000001100000000,
31'b0001100000100000000000000000001,
31'b1000000000001000000000000001100,
31'b1000100100000000010000000010000,
31'b1000000101000001000000010000000,
31'b1001000001000000000000000010100,
31'b1000000000000000000000000001100,
31'b1000000000000010000000000001100,
31'b1000000000000100000000000001100,
31'b1000100000100001000000000000000,
31'b1000000100000000000000101000001,
31'b0110000000000000000011010000000,
31'b0100011000000000010001000000000,
31'b0100000001000001100000000000000,
31'b1000000000010000000000000001100,
31'b1000110010000000000000001000000,
31'b1000000000010100000000000001100,
31'b1000100000110001000000000000000,
31'b1001000100000000000100000000000,
31'b1001000100000010000100000000000,
31'b1001000100000100000100000000000,
31'b1000100000001001000000000000000,
31'b0010001000000000000001000000000,
31'b1000100000000101000000000000000,
31'b1000100000000011000000000000000,
31'b1000100000000001000000000000000,
31'b1001000100010000000100000000000,
31'b0010000000000001000100000000010,
31'b0001000000000010001001000000000,
31'b0001000000000000001001000000000,
31'b1000000000000000001000001000010,
31'b1000100000010101000000000000000,
31'b1000100000010011000000000000000,
31'b1000100000010001000000000000000,
31'b1000000100000101000000010000000,
31'b1001000000000100000000000010100,
31'b1000000100000001000000010000000,
31'b1001000000000000000000000010100,
31'b1000000001000000000000000001100,
31'b1001100000000000000100010000000,
31'b1000000100001001000000010000000,
31'b1001000000001000000000000010100,
31'b0100110010000000000010000000000,
31'b0100000000000101100000000000000,
31'b0100000000000011100000000000000,
31'b0100000000000001100000000000000,
31'b1010000000000000000001011000000,
31'b0100000100000000000010100000001,
31'b0100010000000000000100000100001,
31'b0100000000001001100000000000000,
31'b1001000101000000000100000000000,
31'b0100010010000000100000001000000,
31'b1000100000000000010100000000100,
31'b1001000000100000000000000010100,
31'b1000000000000000010000010010000,
31'b1000100001000101000000000000000,
31'b1000100001000011000000000000000,
31'b1000100001000001000000000000000,
31'b0100100000000000100000000001100,
31'b0100000000000000001010000000010,
31'b0100010000000000001000001001000,
31'b0100000000100001100000000000000,
31'b0010000000000000010000000000110,
31'b0100000100000000110000000010000,
31'b0011000010000000000001100000000,
31'b1100000000000000001000000010001,
31'b0000100000000000000000000000000,
31'b0000100000000010000000000000000,
31'b0000100000000100000000000000000,
31'b0000100000000110000000000000000,
31'b0000100000001000000000000000000,
31'b0000100000001010000000000000000,
31'b0000100000001100000000000000000,
31'b0001000100000001000100000000000,
31'b0000100000010000000000000000000,
31'b0000100000010010000000000000000,
31'b0000100000010100000000000000000,
31'b0000100000010110000000000000000,
31'b0000100000011000000000000000000,
31'b1000001100000000000000001000000,
31'b1010000000000000000100000000010,
31'b1010000000000010000100000000010,
31'b0000100000100000000000000000000,
31'b0000100000100010000000000000000,
31'b0000100000100100000000000000000,
31'b0000000000000001000000000001100,
31'b0000100000101000000000000000000,
31'b0000000101000000000000010000000,
31'b0000100000101100000000000000000,
31'b0000000101000100000000010000000,
31'b0000100000110000000000000000000,
31'b0000000000000000100010001000000,
31'b0000100000110100000000000000000,
31'b0000000000010001000000000001100,
31'b1100000001000000100000000000000,
31'b0000000101010000000000010000000,
31'b1100000001000100100000000000000,
31'b0000000101010100000000010000000,
31'b0000100001000000000000000000000,
31'b0000100001000010000000000000000,
31'b0000100001000100000000000000000,
31'b0000100001000110000000000000000,
31'b0000100001001000000000000000000,
31'b0000000100100000000000010000000,
31'b0000100001001100000000000000000,
31'b0001100000000000000000000011000,
31'b0000100001010000000000000000000,
31'b0100000000000000000000011100000,
31'b0100000000000000010000100000010,
31'b0100000000000100000000011100000,
31'b1100000000100000100000000000000,
31'b0000101000000000100000000100000,
31'b1100000000100100100000000000000,
31'b0001100000010000000000000011000,
31'b0000100001100000000000000000000,
31'b0000000100001000000000010000000,
31'b0000100001100100000000000000000,
31'b0000000100001100000000010000000,
31'b0000000100000010000000010000000,
31'b0000000100000000000000010000000,
31'b0000000000000000010100000001000,
31'b0000000100000100000000010000000,
31'b1100000000001000100000000000000,
31'b0000000100011000000000010000000,
31'b1100000000001100100000000000000,
31'b0010000100000000000010000000101,
31'b1100000000000000100000000000000,
31'b0000000100010000000000010000000,
31'b1100000000000100100000000000000,
31'b0000000100010100000000010000000,
31'b0000100010000000000000000000000,
31'b0000100010000010000000000000000,
31'b0000100010000100000000000000000,
31'b0000100010000110000000000000000,
31'b0000100010001000000000000000000,
31'b0000100010001010000000000000000,
31'b0000100010001100000000000000000,
31'b0001100000000000100000100100000,
31'b0000100010010000000000000000000,
31'b0000100010010010000000000000000,
31'b0000000000000000000010000000110,
31'b0000100000000000101000000001000,
31'b1000000000000000000000000010101,
31'b1000001110000000000000001000000,
31'b0010100000000000000000000110000,
31'b0110000000000000011000000000010,
31'b0000100010100000000000000000000,
31'b0000010000000000001000000000010,
31'b0000100010100100000000000000000,
31'b0000010000000100001000000000010,
31'b0000100010101000000000000000000,
31'b0000010000001000001000000000010,
31'b0000100010101100000000000000000,
31'b1100000001000000001000000001000,
31'b0000100010110000000000000000000,
31'b0000010000010000001000000000010,
31'b0000110000000001000000001000000,
31'b0000110000000011000000001000000,
31'b1100000011000000100000000000000,
31'b0001010100000000000100001000000,
31'b0011011000000000000000000000010,
31'b1110001000000000000000000010000,
31'b0000100011000000000000000000000,
31'b0010010000000000000001010000000,
31'b0000100011000100000000000000000,
31'b0010101000000000100000000010000,
31'b0000100011001000000000000000000,
31'b0010100000000000001000100000000,
31'b0000101000000000001000000101000,
31'b1100000000100000001000000001000,
31'b0101000000000000000001000000100,
31'b0101000000000010000001000000100,
31'b0001101000000000000000100000000,
31'b1001000000000000000000000001101,
31'b1100000010100000100000000000000,
31'b0010100000010000001000100000000,
31'b0010100001000000000000000110000,
31'b1100000000000000000000001000110,
31'b0000100011100000000000000000000,
31'b0000010001000000001000000000010,
31'b0000101000000000000100001000001,
31'b1100000000001000001000000001000,
31'b0000000000000000001001000000001,
31'b0000000110000000000000010000000,
31'b0000000010000000010100000001000,
31'b1100000000000000001000000001000,
31'b1100000010001000100000000000000,
31'b0000010001010000001000000000010,
31'b0011000000000001000000000100100,
31'b1101000000000000000000100100000,
31'b1100000010000000100000000000000,
31'b0000000110010000000000010000000,
31'b1100000010000100100000000000000,
31'b1000000100000000000100000000001,
31'b0000100100000000000000000000000,
31'b0000100100000010000000000000000,
31'b0000100100000100000000000000000,
31'b0001000000001001000100000000000,
31'b0000100100001000000000000000000,
31'b0000000001100000000000010000000,
31'b0001000000000011000100000000000,
31'b0001000000000001000100000000000,
31'b0000100100010000000000000000000,
31'b1000001000001000000000001000000,
31'b0001001000000000000001000000010,
31'b1000100000000000001101000000000,
31'b1000001000000010000000001000000,
31'b1000001000000000000000001000000,
31'b1010000100000000000100000000010,
31'b1000001000000100000000001000000,
31'b0000100100100000000000000000000,
31'b0000000001001000000000010000000,
31'b0001000000000000000000010011000,
31'b0000000100000001000000000001100,
31'b0000000001000010000000010000000,
31'b0000000001000000000000010000000,
31'b0000100000000001010000000010000,
31'b0000000001000100000000010000000,
31'b0000100100110000000000000000000,
31'b0000000100000000100010001000000,
31'b0001001000100000000001000000010,
31'b0010000001000000000010000000101,
31'b0100100000000000000000001100000,
31'b0000000001010000000000010000000,
31'b0100100000000100000000001100000,
31'b0000000001010100000000010000000,
31'b0000100101000000000000000000000,
31'b0000000000101000000000010000000,
31'b0001000000000000010000000000100,
31'b0001000000000010010000000000100,
31'b0000000000100010000000010000000,
31'b0000000000100000000000010000000,
31'b0001000000001000010000000000100,
31'b0000000000100100000000010000000,
31'b0100001000000000000010000000000,
31'b0100001000000010000010000000000,
31'b0100001000000100000010000000000,
31'b0110010000000000010000010000000,
31'b0100001000001000000010000000000,
31'b0000000000110000000000010000000,
31'b0100001000001100000010000000000,
31'b0001011000000000000000000000001,
31'b0000000000001010000000010000000,
31'b0000000000001000000000010000000,
31'b0001000000100000010000000000100,
31'b0000000000001100000000010000000,
31'b0000000000000010000000010000000,
31'b0000000000000000000000010000000,
31'b0000000000000110000000010000000,
31'b0000000000000100000000010000000,
31'b0100001000100000000010000000000,
31'b0000000000011000000000010000000,
31'b0100001000100100000010000000000,
31'b0010000000000000000010000000101,
31'b0000000000010010000000010000000,
31'b0000000000010000000000010000000,
31'b0100000000000000011000000000001,
31'b0000000000010100000000010000000,
31'b0000100110000000000000000000000,
31'b0000100110000010000000000000000,
31'b0101000000000000000010100000000,
31'b0101000000000010000010100000000,
31'b0000100110001000000000000000000,
31'b0000010000000000000000100000001,
31'b0101000000001000000010100000000,
31'b0001000010000001000100000000000,
31'b0000100110010000000000000000000,
31'b1000100000000000010000000001001,
31'b0100100000000000010001000000000,
31'b0110000000000000100010000010000,
31'b1000001010000010000000001000000,
31'b1000001010000000000000001000000,
31'b0100100000001000010001000000000,
31'b1000001010000100000000001000000,
31'b0010000000000000001000110000000,
31'b0000010100000000001000000000010,
31'b0110100000000000000000001010000,
31'b1000011000001001000000000000000,
31'b0010110000000000000001000000000,
31'b0000000011000000000000010000000,
31'b1000011000000011000000000000000,
31'b1000011000000001000000000000000,
31'b0010100000000001010000000100000,
31'b0001010000001000000100001000000,
31'b1000010000000000000101000000010,
31'b1000001000000000010001000100000,
31'b0100100010000000000000001100000,
31'b0001010000000000000100001000000,
31'b1000001000000000100000000000110,
31'b1000000001000000000100000000001,
31'b0000000000000000000001100000010,
31'b0000000010101000000000010000000,
31'b0001000010000000010000000000100,
31'b1001000000001000000000101000000,
31'b0000000010100010000000010000000,
31'b0000000010100000000000010000000,
31'b1001000000000010000000101000000,
31'b1001000000000000000000101000000,
31'b0100001010000000000010000000000,
31'b0100001010000010000010000000000,
31'b0100100001000000010001000000000,
31'b1000000000101000000100000000001,
31'b0100001010001000000010000000000,
31'b0000001000000001000100100000000,
31'b1010000000000000100000001010000,
31'b1000000000100000000100000000001,
31'b0000000010001010000000010000000,
31'b0000000010001000000000010000000,
31'b1000000000001000110001000000000,
31'b1000000000000000000000000100110,
31'b0000000010000010000000010000000,
31'b0000000010000000000000010000000,
31'b1000000000000000110001000000000,
31'b0000000010000100000000010000000,
31'b0100001010100000000010000000000,
31'b0000000010011000000000010000000,
31'b1000010000000001100000000100000,
31'b1000000000001000000100000000001,
31'b0100000000000000000101000001000,
31'b0000000010010000000000010000000,
31'b1000000000000010000100000000001,
31'b1000000000000000000100000000001,
31'b0000101000000000000000000000000,
31'b0000101000000010000000000000000,
31'b0000101000000100000000000000000,
31'b1010000000000001000001000000000,
31'b0000101000001000000000000000000,
31'b1000000100010000000000001000000,
31'b0000101000001100000000000000000,
31'b1010000000001001000001000000000,
31'b0000101000010000000000000000000,
31'b1000000100001000000000001000000,
31'b0001000100000000000001000000010,
31'b1010000000010001000001000000000,
31'b1000000100000010000000001000000,
31'b1000000100000000000000001000000,
31'b1010001000000000000100000000010,
31'b1000000100000100000000001000000,
31'b0000101000100000000000000000000,
31'b1100000000000000000000000100000,
31'b0000101000100100000000000000000,
31'b1100000000000100000000000100000,
31'b0000101000101000000000000000000,
31'b1100000000001000000000000100000,
31'b0000101000101100000000000000000,
31'b1100000000001100000000000100000,
31'b0000101000110000000000000000000,
31'b1100000000010000000000000100000,
31'b0001110000000000000000010000001,
31'b1100000000010100000000000100000,
31'b1100001001000000100000000000000,
31'b1000000100100000000000001000000,
31'b0011010010000000000000000000010,
31'b1110000010000000000000000010000,
31'b0000101001000000000000000000000,
31'b1000000000000000100010010000000,
31'b0000101001000100000000000000000,
31'b1010000001000001000001000000000,
31'b0000101001001000000000000000000,
31'b0000100000010000100000000100000,
31'b0000101001001100000000000000000,
31'b0001101000000000000000000011000,
31'b0100000100000000000010000000000,
31'b0100000100000010000010000000000,
31'b0100000100000100000010000000000,
31'b0100010000000000000100100100000,
31'b0100000100001000000010000000000,
31'b0000100000000000100000000100000,
31'b0100000100001100000010000000000,
31'b0001010100000000000000000000001,
31'b0000101001100000000000000000000,
31'b1100000001000000000000000100000,
31'b0000101001100100000000000000000,
31'b1100000001000100000000000100000,
31'b0000000000000000000010001100000,
31'b0000001100000000000000010000000,
31'b0000001000000000010100000001000,
31'b0000010000000000000000000101010,
31'b1000100000000000000000011000000,
31'b1100000001010000000000000100000,
31'b1100000000000000001000100010000,
31'b0011000010000000000001000000001,
31'b1100001000000000100000000000000,
31'b0000100000100000100000000100000,
31'b1100001000000100100000000000000,
31'b0001100000000000000001010000010,
31'b0000101010000000000000000000000,
31'b1000010000000000010000000010000,
31'b0000101010000100000000000000000,
31'b1010000010000001000001000000000,
31'b0000101010001000000000000000000,
31'b1000010000001000010000000010000,
31'b0000101010001100000000000000000,
31'b1100000000000000010001001000000,
31'b0000101010010000000000000000000,
31'b1000010000010000010000000010000,
31'b0001100001000000000000100000000,
31'b0001100001000010000000100000000,
31'b1000001000000000000000000010101,
31'b1000000110000000000000001000000,
31'b0011010000100000000000000000010,
31'b1110000000100000000000000010000,
31'b0000101010100000000000000000000,
31'b1100000010000000000000000100000,
31'b0000101010100100000000000000000,
31'b1100000010000100000000000100000,
31'b0000101010101000000000000000000,
31'b1100000010001000000000000100000,
31'b1101000000000000100000100000000,
31'b1000010100000001000000000000000,
31'b0000101010110000000000000000000,
31'b1100000010010000000000000100000,
31'b0011010000001000000000000000010,
31'b1110000000001000000000000010000,
31'b0011010000000100000000000000010,
31'b1110000000000100000000000010000,
31'b0011010000000000000000000000010,
31'b1110000000000000000000000010000,
31'b0000101011000000000000000000000,
31'b1000010001000000010000000010000,
31'b0000000000000000010011000000000,
31'b0010100000000000100000000010000,
31'b0000101011001000000000000000000,
31'b0010101000000000001000100000000,
31'b0000100000000000001000000101000,
31'b0110000000000000001001000000100,
31'b0100000110000000000010000000000,
31'b0101000000000001000000000100001,
31'b0001100000000000000000100000000,
31'b0001100000000010000000100000000,
31'b0101010000000000100100000000000,
31'b0000100010000000100000000100000,
31'b0001100000001000000000100000000,
31'b0001100000001010000000100000000,
31'b0000101011100000000000000000000,
31'b1100000011000000000000000100000,
31'b0000100000000000000100001000001,
31'b0011000000010000000001000000001,
31'b0000001000000000001001000000001,
31'b0000001110000000000000010000000,
31'b0000100000100000001000000101000,
31'b1100001000000000001000000001000,
31'b1111000000000000000000000001000,
31'b0011000000000100000001000000001,
31'b0010000000000000000010001010000,
31'b0011000000000000000001000000001,
31'b1100001010000000100000000000000,
31'b0000100010100000100000000100000,
31'b0011010001000000000000000000010,
31'b1110000001000000000000000010000,
31'b0000101100000000000000000000000,
31'b1000000000011000000000001000000,
31'b0001000000010000000001000000010,
31'b1010000100000001000001000000000,
31'b1000000000010010000000001000000,
31'b1000000000010000000000001000000,
31'b1000100000000001001000000000010,
31'b1000000000010100000000001000000,
31'b0100000001000000000010000000000,
31'b1000000000001000000000001000000,
31'b0001000000000000000001000000010,
31'b1000000000001100000000001000000,
31'b1000000000000010000000001000000,
31'b1000000000000000000000001000000,
31'b1000000000000110000000001000000,
31'b1000000000000100000000001000000,
31'b0000101100100000000000000000000,
31'b1100000100000000000000000100000,
31'b0001001000000000000000010011000,
31'b1100000100000100000000000100000,
31'b1000100000000000100010000000000,
31'b0000001001000000000000010000000,
31'b1000100000000100100010000000000,
31'b1000010010000001000000000000000,
31'b0000000000000000100000010100000,
31'b1000000000101000000000001000000,
31'b0001000000100000000001000000010,
31'b1000000010000000010001000100000,
31'b1000000000100010000000001000000,
31'b1000000000100000000000001000000,
31'b1000000010000000100000000000110,
31'b1000000000100100000000001000000,
31'b0100000000010000000010000000000,
31'b0100000000010010000010000000000,
31'b0100000000010100000010000000000,
31'b0100010000100000001000000000100,
31'b0100000000011000000010000000000,
31'b0000001000100000000000010000000,
31'b0110000000000000000000010000101,
31'b0001010000010000000000000000001,
31'b0100000000000000000010000000000,
31'b0100000000000010000010000000000,
31'b0100000000000100000010000000000,
31'b0100000000000110000010000000000,
31'b0100000000001000000010000000000,
31'b1000000001000000000000001000000,
31'b0100000000001100000010000000000,
31'b0001010000000000000000000000001,
31'b0100000000110000000010000000000,
31'b0000001000001000000000010000000,
31'b0100010000000010001000000000100,
31'b0100010000000000001000000000100,
31'b0000001000000010000000010000000,
31'b0000001000000000000000010000000,
31'b0010010000000000010010000000000,
31'b0000001000000100000000010000000,
31'b0100000000100000000010000000000,
31'b0100000000100010000010000000000,
31'b0100000000100100000010000000000,
31'b0100010000010000001000000000100,
31'b0100000000101000000010000000000,
31'b0000001000010000000000010000000,
31'b0100001000000000011000000000001,
31'b0001010000100000000000000000001,
31'b0000101110000000000000000000000,
31'b1000010100000000010000000010000,
31'b0101001000000000000010100000000,
31'b1010000000000000000000001110000,
31'b1000110000000000000000000001100,
31'b1000000010010000000000001000000,
31'b1000010000100011000000000000000,
31'b1000010000100001000000000000000,
31'b0000000000000000010000100000100,
31'b1000000010001000000000001000000,
31'b0001000010000000000001000000010,
31'b1000000010001100000000001000000,
31'b1000000010000010000000001000000,
31'b1000000010000000000000001000000,
31'b1000000010000110000000001000000,
31'b1000000010000100000000001000000,
31'b0010100000000000100100000000100,
31'b1100000110000000000000000100000,
31'b1000010000001011000000000000000,
31'b1000010000001001000000000000000,
31'b1000100010000000100010000000000,
31'b1000010000000101000000000000000,
31'b1000010000000011000000000000000,
31'b1000010000000001000000000000000,
31'b0000000010000000100000010100000,
31'b1000000010101000000000001000000,
31'b1000000000001000100000000000110,
31'b1000000000000000010001000100000,
31'b1000000010100010000000001000000,
31'b1000000010100000000000001000000,
31'b1000000000000000100000000000110,
31'b0001000000000000000000110000000,
31'b0100000010010000000010000000000,
31'b0100000010010010000010000000000,
31'b0100100000000000000000000000110,
31'b0100100000000010000000000000110,
31'b0100000010011000000010000000000,
31'b0000001010100000000000010000000,
31'b0110000000000000000010000110000,
31'b1001001000000000000000101000000,
31'b0100000010000000000010000000000,
31'b0100000010000010000010000000000,
31'b0100000010000100000010000000000,
31'b0100110000000001100000000000000,
31'b0100000010001000000010000000000,
31'b0000000000000001000100100000000,
31'b0100100000000000000100000100001,
31'b0001010010000000000000000000001,
31'b0100000010110000000010000000000,
31'b0100000000000001000000000001010,
31'b1000010000000000010100000000100,
31'b1000010001001001000000000000000,
31'b0000001010000010000000010000000,
31'b0000001010000000000000010000000,
31'b1000010001000011000000000000000,
31'b1000010001000001000000000000000,
31'b0100000010100000000010000000000,
31'b0100000010100010000010000000000,
31'b0100100000000000001000001001000,
31'b1000001000001000000100000000001,
31'b0100001000000000000101000001000,
31'b0000001010010000000000010000000,
31'b1000001000000010000100000000001,
31'b1000001000000000000100000000001,
31'b0000110000000000000000000000000,
31'b0000110000000010000000000000000,
31'b0000110000000100000000000000000,
31'b0000110000000110000000000000000,
31'b0000110000001000000000000000000,
31'b0000110000001010000000000000000,
31'b0100000000000000100100100000000,
31'b0101100000000000000010000000001,
31'b0000110000010000000000000000000,
31'b0000110000010010000000000000000,
31'b0000110000010100000000000000000,
31'b0000110000010110000000000000000,
31'b1000000000000000010000100001000,
31'b1000011100000000000000001000000,
31'b1010010000000000000100000000010,
31'b1010001000000000010000000100000,
31'b0000110000100000000000000000000,
31'b0000000010000000001000000000010,
31'b0000110000100100000000000000000,
31'b0000010000000001000000000001100,
31'b0010000001000000000000100000010,
31'b0000010101000000000000010000000,
31'b0110100000010000010000000000000,
31'b1000001110000001000000000000000,
31'b0000110000110000000000000000000,
31'b0000010000000000100010001000000,
31'b0000000000000000100000000001010,
31'b0000100000000000001010000000100,
31'b1100010001000000100000000000000,
31'b0001000110000000000100001000000,
31'b0110100000000000010000000000000,
31'b0110100000000010010000000000000,
31'b0000110001000000000000000000000,
31'b0010000010000000000001010000000,
31'b1010000000000000110000000000000,
31'b1010000000000010110000000000000,
31'b0010000000100000000000100000010,
31'b0000100000000000000001000000011,
31'b1100100000000000000000000001010,
31'b0001110000000000000000000011000,
31'b0110000000000000000100000001000,
31'b0110000000000010000100000001000,
31'b1010000000010000110000000000000,
31'b1010000000000000000101000000001,
31'b1100010000100000100000000000000,
31'b0001001100000100000000000000001,
31'b0001001100000010000000000000001,
31'b0001001100000000000000000000001,
31'b0010000000001000000000100000010,
31'b0000010100001000000000010000000,
31'b1010000000100000110000000000000,
31'b0100001100000000001000000000100,
31'b0010000000000000000000100000010,
31'b0000010100000000000000010000000,
31'b0010000000000100000000100000010,
31'b0000010100000100000000010000000,
31'b1100010000001000100000000000000,
31'b0001000100000000011010000000000,
31'b1000100000000000000100100000000,
31'b1001000000000000100010000000001,
31'b1100010000000000100000000000000,
31'b0001000000000000100000000010010,
31'b1100010000000100100000000000000,
31'b0001001100100000000000000000001,
31'b0000110010000000000000000000000,
31'b0000000000100000001000000000010,
31'b0000110010000100000000000000000,
31'b0000000000000001100010000000000,
31'b0000110010001000000000000000000,
31'b0000000100000000000000100000001,
31'b0100100100000001000000000100000,
31'b0000000100000100000000100000001,
31'b0000110010010000000000000000000,
31'b0000000000000000000000001001100,
31'b0000100000100001000000001000000,
31'b0000000000010001100010000000000,
31'b1000010000000000000000000010101,
31'b0000000100010000000000100000001,
31'b0011001000100000000000000000010,
31'b0000000101000001000000011000000,
31'b0000000000000010001000000000010,
31'b0000000000000000001000000000010,
31'b0000100000010001000000001000000,
31'b0000000000000100001000000000010,
31'b0010100100000000000001000000000,
31'b0000000000001000001000000000010,
31'b1001000000000000001001001000000,
31'b1000001100000001000000000000000,
31'b0000100000000101000000001000000,
31'b0000000000010000001000000000010,
31'b0000100000000001000000001000000,
31'b0000100000000011000000001000000,
31'b0011001000000100000000000000010,
31'b0001000100000000000100001000000,
31'b0011001000000000000000000000010,
31'b1010100000000000001100000000000,
31'b0010000000000010000001010000000,
31'b0010000000000000000001010000000,
31'b1010000010000000110000000000000,
31'b0010000000000100000001010000000,
31'b0010000010100000000000100000010,
31'b0010000000001000000001010000000,
31'b1100000000000001100000001000000,
31'b0010000000001100000001010000000,
31'b0110000010000000000100000001000,
31'b0010000000010000000001010000000,
31'b0001111000000000000000100000000,
31'b0010000100000000100000000001001,
31'b1100000000000000000010000001100,
31'b0010000000011000000001010000000,
31'b0001000000000000000000001010100,
31'b0000000100000001000000011000000,
31'b0000100000000000000000110000001,
31'b0000000001000000001000000000010,
31'b0100000000000011000000010100000,
31'b0100000000000001000000010100000,
31'b0010000010000000000000100000010,
31'b0000010110000000000000010000000,
31'b0011000000000000010001000000100,
31'b1100010000000000001000000001000,
31'b0000100001000101000000001000000,
31'b0000000001010000001000000000010,
31'b0000100001000001000000001000000,
31'b0100100000000000011000100000000,
31'b1100010010000000100000000000000,
31'b0001000101000000000100001000000,
31'b0011001001000000000000000000010,
31'b1100100000000001000010000000000,
31'b0000110100000000000000000000000,
31'b0000110100000010000000000000000,
31'b0001000000000000100000000100001,
31'b0001010000001001000100000000000,
31'b0000110100001000000000000000000,
31'b0000000010000000000000100000001,
31'b0100100010000001000000000100000,
31'b0001010000000001000100000000000,
31'b0000110100010000000000000000000,
31'b1000100000000000000000100010100,
31'b0001011000000000000001000000010,
31'b1100001000000000000001000010000,
31'b1000011000000010000000001000000,
31'b1000011000000000000000001000000,
31'b1000001000000000000010000001010,
31'b1000000000000000000100110000000,
31'b0000110100100000000000000000000,
31'b0000010001001000000000010000000,
31'b0001010000000000000000010011000,
31'b1100000000000000000000010001010,
31'b0010100010000000000001000000000,
31'b0000010001000000000000010000000,
31'b1000001010000011000000000000000,
31'b1000001010000001000000000000000,
31'b0000110100110000000000000000000,
31'b0001000010001000000100001000000,
31'b0000100000000000000001000110000,
31'b0110000000000000000000000011100,
31'b0111000001000000000000000000100,
31'b0001000010000000000100001000000,
31'b0110100100000000010000000000000,
31'b1000001010010001000000000000000,
31'b0010000000000000001000000000001,
31'b0010000000000010001000000000001,
31'b0010000000000100001000000000001,
31'b0110000000010000010000010000000,
31'b0010000000001000001000000000001,
31'b0000010000100000000000010000000,
31'b0010001000100000010010000000000,
31'b0001001000010000000000000000001,
31'b0100011000000000000010000000000,
31'b0110000000000100010000010000000,
31'b0110000000000010010000010000000,
31'b0110000000000000010000010000000,
31'b0111000000100000000000000000100,
31'b0001001000000100000000000000001,
31'b0001001000000010000000000000001,
31'b0001001000000000000000000000001,
31'b0010000000100000001000000000001,
31'b0000010000001000000000010000000,
31'b0101000000000000000010010000001,
31'b0100001000000000001000000000100,
31'b0000010000000010000000010000000,
31'b0000010000000000000000010000000,
31'b0010001000000000010010000000000,
31'b0000010000000100000000010000000,
31'b0111000000001000000000000000100,
31'b0001000000000000011010000000000,
31'b1000100100000000000100100000000,
31'b0110000000100000010000010000000,
31'b0111000000000000000000000000100,
31'b0000010000010000000000010000000,
31'b0111000000000100000000000000100,
31'b0001001000100000000000000000001,
31'b0000110110000000000000000000000,
31'b0000000000001000000000100000001,
31'b0101010000000000000010100000000,
31'b0000000100000001100010000000000,
31'b0000000000000010000000100000001,
31'b0000000000000000000000100000001,
31'b0100100000000001000000000100000,
31'b0000000000000100000000100000001,
31'b0000110110010000000000000000000,
31'b0000000100000000000000001001100,
31'b1100000000000001000010010000000,
31'b0010000001000000100000000001001,
31'b0000100000000000010000001010000,
31'b0000000000010000000000100000001,
31'b0100100000010001000000000100000,
31'b0000000001000001000000011000000,
31'b0010100000001000000001000000000,
31'b0000000100000000001000000000010,
31'b1000001000001011000000000000000,
31'b1000001000001001000000000000000,
31'b0010100000000000000001000000000,
31'b0000000000100000000000100000001,
31'b1000001000000011000000000000000,
31'b1000001000000001000000000000000,
31'b1011000000000001001000000000000,
31'b0001000000001000000100001000000,
31'b1000000000000000000101000000010,
31'b1000001000011001000000000000000,
31'b0010100000010000000001000000000,
31'b0001000000000000000100001000000,
31'b1000001000010011000000000000000,
31'b1000001000010001000000000000000,
31'b0010000010000000001000000000001,
31'b0010000100000000000001010000000,
31'b0010000010000100001000000000001,
31'b0010000100000100000001010000000,
31'b0000100000000000001000010000010,
31'b0000000001000000000000100000001,
31'b0100100001000001000000000100000,
31'b0000000001000100000000100000001,
31'b1110000000000000100001000000000,
31'b0010000100010000000001010000000,
31'b1010000000000000001100010000000,
31'b0010000000000000100000000001001,
31'b0000100001000000010000001010000,
31'b0000000001010000000000100000001,
31'b0000000000000011000000011000000,
31'b0000000000000001000000011000000,
31'b0010100001001000000001000000000,
31'b0000010010001000000000010000000,
31'b1000001000000000010100000000100,
31'b1000010000000000000000000100110,
31'b0010100001000000000001000000000,
31'b0000010010000000000000010000000,
31'b1000010000000000110001000000000,
31'b1000001001000001000000000000000,
31'b1101000000000000000110000000000,
31'b0001000010000000011010000000000,
31'b1000000000000001100000000100000,
31'b1000010000001000000100000000001,
31'b0111000010000000000000000000100,
31'b0001000001000000000100001000000,
31'b1000010000000010000100000000001,
31'b1000010000000000000100000000001,
31'b0000111000000000000000000000000,
31'b1000000010000000010000000010000,
31'b0000111000000100000000000000000,
31'b1010010000000001000001000000000,
31'b0000111000001000000000000000000,
31'b1000010100010000000000001000000,
31'b0100100000000000001000010000100,
31'b1010000000010000010000000100000,
31'b0000111000010000000000000000000,
31'b1000010100001000000000001000000,
31'b0001100000100000000000010000001,
31'b1100000100000000000001000010000,
31'b1000010100000010000000001000000,
31'b1000010100000000000000001000000,
31'b1010000000000010010000000100000,
31'b1010000000000000010000000100000,
31'b0001000000000000000000000110010,
31'b1100010000000000000000000100000,
31'b0001100000010000000000010000001,
31'b1100010000000100000000000100000,
31'b0011100000000000000010000000100,
31'b1100010000001000000000000100000,
31'b1001000000000000000010000100001,
31'b1000000110000001000000000000000,
31'b0001100000000100000000010000001,
31'b1100010000010000000000000100000,
31'b0001100000000000000000010000001,
31'b0001100000000010000000010000001,
31'b0011000010000100000000000000010,
31'b1100000000000001010001000000000,
31'b0011000010000000000000000000010,
31'b1010000000100000010000000100000,
31'b0010000000000001000010000010000,
31'b1000010000000000100010010000000,
31'b1010001000000000110000000000000,
31'b0100000100100000001000000000100,
31'b0010001000100000000000100000010,
31'b0001000100010100000000000000001,
31'b1010000000000001000000000000011,
31'b0001000100010000000000000000001,
31'b0100010100000000000010000000000,
31'b0100010100000010000010000000000,
31'b0100010100000100000010000000000,
31'b0100000000000000000100100100000,
31'b0101000010000000100100000000000,
31'b0001000100000100000000000000001,
31'b0001000100000010000000000000001,
31'b0001000100000000000000000000001,
31'b0010001000001000000000100000010,
31'b1100010001000000000000000100000,
31'b0100000100000010001000000000100,
31'b0100000100000000001000000000100,
31'b0010001000000000000000100000010,
31'b0000011100000000000000010000000,
31'b0010000100000000010010000000000,
31'b0000000000000000000000000101010,
31'b1100000000000000000101000000100,
31'b0010000010000000000000000011010,
31'b1000101000000000000100100000000,
31'b0001000000000000001000100000010,
31'b1100011000000000100000000000000,
31'b0001001000000000100000000010010,
31'b0011000011000000000000000000010,
31'b0001000100100000000000000000001,
31'b1000000000000010010000000010000,
31'b1000000000000000010000000010000,
31'b1000100001000001000000010000000,
31'b1000000000000100010000000010000,
31'b1000100100000000000000000001100,
31'b1000000000001000010000000010000,
31'b1001000001000000010000000001000,
31'b1000000100100001000000000000000,
31'b1000100000000000000000101000001,
31'b1000000000010000010000000010000,
31'b0011000000101000000000000000010,
31'b1100000000000001000000001100000,
31'b0101000001000000100100000000000,
31'b1000010110000000000000001000000,
31'b0011000000100000000000000000010,
31'b1010000010000000010000000100000,
31'b1001100000000000000100000000000,
31'b0000001000000000001000000000010,
31'b1001100000000100000100000000000,
31'b1000000100001001000000000000000,
31'b1001100000001000000100000000000,
31'b1000000100000101000000000000000,
31'b1000000100000011000000000000000,
31'b1000000100000001000000000000000,
31'b1010000000000010000001001000000,
31'b1010000000000000000001001000000,
31'b0011000000001000000000000000010,
31'b1010000000000100000001001000000,
31'b0011000000000100000000000000010,
31'b1010000000001000000001001000000,
31'b0011000000000000000000000000010,
31'b1000000100010001000000000000000,
31'b1000100000000101000000010000000,
31'b1000000001000000010000000010000,
31'b1000100000000001000000010000000,
31'b1000100000000011000000010000000,
31'b1001000000000100010000000001000,
31'b1001000100000000000100010000000,
31'b1001000000000000010000000001000,
31'b1001000000000010010000000001000,
31'b0101000000001000100100000000000,
31'b1000000001010000010000000010000,
31'b0001110000000000000000100000000,
31'b0100100100000001100000000000000,
31'b0101000000000000100100000000000,
31'b0101000000000010100100000000000,
31'b0000000000000001000010000100000,
31'b0001000110000000000000000000001,
31'b1001100001000000000100000000000,
31'b1000000000000000000000010001100,
31'b1000100000100001000000010000000,
31'b1000000101001001000000000000000,
31'b0110000000010000000011000000000,
31'b1000000101000101000000000000000,
31'b1001000000100000010000000001000,
31'b1000000101000001000000000000000,
31'b0110000000001000000011000000000,
31'b0010000000000000000000000011010,
31'b0011000001001000000000000000010,
31'b0011010000000000000001000000001,
31'b0110000000000000000011000000000,
31'b0110000000000010000011000000000,
31'b0011000001000000000000000000010,
31'b1010000000000000000010000001001,
31'b0000111100000000000000000000000,
31'b1000010000011000000000001000000,
31'b0001010000010000000001000000010,
31'b1100000000010000000001000010000,
31'b1000100010000000000000000001100,
31'b1000010000010000000000001000000,
31'b1000000010100011000000000000000,
31'b1000000010100001000000000000000,
31'b0000000000000000000000000011001,
31'b1000010000001000000000001000000,
31'b0001010000000000000001000000010,
31'b1100000000000000000001000010000,
31'b1000010000000010000000001000000,
31'b1000010000000000000000001000000,
31'b1000000000000000000010000001010,
31'b0001000001000000000000000000001,
31'b0001100000000000100001000001000,
31'b1100010100000000000000000100000,
31'b1100000000000000000110100000000,
31'b1000000010001001000000000000000,
31'b1000110000000000100010000000000,
31'b1000000010000101000000000000000,
31'b1000000010000011000000000000000,
31'b1000000010000001000000000000000,
31'b0000010000000000100000010100000,
31'b1010000000000001000000000110000,
31'b0001100100000000000000010000001,
31'b1100000000100000000001000010000,
31'b1000010000100010000000001000000,
31'b1000010000100000000000001000000,
31'b1000000010010011000000000000000,
31'b1000000010010001000000000000000,
31'b0100010000010000000010000000000,
31'b0100010000010010000010000000000,
31'b0100010000010100000010000000000,
31'b0100000000100000001000000000100,
31'b0101000000000000011000010000000,
31'b0001000000010100000000000000001,
31'b0010000000100000010010000000000,
31'b0001000000010000000000000000001,
31'b0100010000000000000010000000000,
31'b0100010000000010000010000000000,
31'b0100010000000100000010000000000,
31'b0001000000001000000000000000001,
31'b0100010000001000000010000000000,
31'b0001000000000100000000000000001,
31'b0001000000000010000000000000001,
31'b0001000000000000000000000000001,
31'b0100010000110000000010000000000,
31'b0100000000000100001000000000100,
31'b0100000000000010001000000000100,
31'b0100000000000000001000000000100,
31'b0010000000000100010010000000000,
31'b0000011000000000000000010000000,
31'b0010000000000000010010000000000,
31'b0000000000000000000100101000000,
31'b0100010000100000000010000000000,
31'b0100010000100010000010000000000,
31'b0100010000100100000010000000000,
31'b0100000000010000001000000000100,
31'b0111001000000000000000000000100,
31'b0001000000100100000000000000001,
31'b0010000000010000010010000000000,
31'b0001000000100000000000000000001,
31'b1000100000001000000000000001100,
31'b1000000100000000010000000010000,
31'b1000000000101011000000000000000,
31'b1000000000101001000000000000000,
31'b1000100000000000000000000001100,
31'b0000001000000000000000100000001,
31'b1000000000100011000000000000000,
31'b1000000000100001000000000000000,
31'b0000010000000000010000100000100,
31'b1000010010001000000000001000000,
31'b0011000000000000001000100000001,
31'b1100000010000000000001000010000,
31'b1000100000010000000000000001100,
31'b1000010010000000000000001000000,
31'b1000000010000000000010000001010,
31'b1000000000110001000000000000000,
31'b1001100100000000000100000000000,
31'b1000000000001101000000000000000,
31'b1000000000001011000000000000000,
31'b1000000000001001000000000000000,
31'b1000000000000111000000000000000,
31'b1000000000000101000000000000000,
31'b1000000000000011000000000000000,
31'b1000000000000001000000000000000,
31'b0100000001000000100000000001100,
31'b1010000100000000000001001000000,
31'b1000001000000000000101000000010,
31'b1000000000011001000000000000000,
31'b1000100000000000001000001000010,
31'b1000000000010101000000000000000,
31'b1000000000010011000000000000000,
31'b1000000000010001000000000000000,
31'b0100010010010000000010000000000,
31'b1001000000001000000100010000000,
31'b1000100100000001000000010000000,
31'b1001100000000000000000000010100,
31'b1001000000000010000100010000000,
31'b1001000000000000000100010000000,
31'b1001000100000000010000000001000,
31'b1000000001100001000000000000000,
31'b0100010010000000000010000000000,
31'b0100100000000101100000000000000,
31'b0100100000000011100000000000000,
31'b0100100000000001100000000000000,
31'b0101000100000000100100000000000,
31'b0001000010000100000000000000001,
31'b0001000010000010000000000000001,
31'b0001000010000000000000000000001,
31'b1001000000000001000000000011000,
31'b1000000100000000000000010001100,
31'b1000000000000000010100000000100,
31'b1000000001001001000000000000000,
31'b1000100000000000010000010010000,
31'b1000000001000101000000000000000,
31'b1000000001000011000000000000000,
31'b1000000001000001000000000000000,
31'b0100000000000000100000000001100,
31'b0100100000000000001010000000010,
31'b1000001000000001100000000100000,
31'b1000000001011001000000000000000,
31'b0110000100000000000011000000000,
31'b1000000001010101000000000000000,
31'b1000000001010011000000000000000,
31'b1000000001010001000000000000000,
31'b0001000000000000000000000000000,
31'b0001000000000010000000000000000,
31'b0001000000000100000000000000000,
31'b0001000000000110000000000000000,
31'b0001000000001000000000000000000,
31'b0001000000001010000000000000000,
31'b0001000000001100000000000000000,
31'b0000000001000000000000000011000,
31'b0001000000010000000000000000000,
31'b0001000000010010000000000000000,
31'b0001000000010100000000000000000,
31'b0010001000001000001000000000000,
31'b0001000000011000000000000000000,
31'b0010001000000100001000000000000,
31'b0010001000000010001000000000000,
31'b0010001000000000001000000000000,
31'b0001000000100000000000000000000,
31'b0001000000100010000000000000000,
31'b0001000000100100000000000000000,
31'b0001000000100110000000000000000,
31'b0001000000101000000000000000000,
31'b0001000000101010000000000000000,
31'b0001000000101100000000000000000,
31'b0000000000000000010000010000100,
31'b0001000000110000000000000000000,
31'b0010000000000000010010000000001,
31'b0001000000110100000000000000000,
31'b0010001000101000001000000000000,
31'b0100000000000000001000000000101,
31'b0101001000000000000010010000000,
31'b0111010000000000010000000000000,
31'b0010001000100000001000000000000,
31'b0001000001000000000000000000000,
31'b0001000001000010000000000000000,
31'b0001000001000100000000000000000,
31'b0000000000001000000000000011000,
31'b0001000001001000000000000000000,
31'b0000000000000100000000000011000,
31'b0000000000000010000000000011000,
31'b0000000000000000000000000011000,
31'b0001000001010000000000000000000,
31'b0010000010000000000000000101000,
31'b0000001010000000000000100000000,
31'b0000001010000010000000100000000,
31'b0001000001011000000000000000000,
31'b0001001000000000100000000100000,
31'b0000001010001000000000100000000,
31'b0000000000010000000000000011000,
31'b0001000001100000000000000000000,
31'b0001000001100010000000000000000,
31'b0000000000000001000100010000000,
31'b0000000000101000000000000011000,
31'b0001000001101000000000000000000,
31'b0001100100000000000000010000000,
31'b0000000000100010000000000011000,
31'b0000000000100000000000000011000,
31'b1000000010000001000000000000001,
31'b1001000100000000000010000100000,
31'b0000001010100000000000100000000,
31'b0100000010000001000001000001000,
31'b1101100000000000100000000000000,
31'b0001100100010000000000010000000,
31'b0000001010101000000000100000000,
31'b0000001000000000000001010000010,
31'b0001000010000000000000000000000,
31'b0001000010000010000000000000000,
31'b0001000010000100000000000000000,
31'b0001000010000110000000000000000,
31'b0001000010001000000000000000000,
31'b0001000010001010000000000000000,
31'b0001000010001100000000000000000,
31'b0000000000000000100000100100000,
31'b0001000010010000000000000000000,
31'b0010000001000000000000000101000,
31'b0000001001000000000000100000000,
31'b0001000000000000101000000001000,
31'b0001000010011000000000000000000,
31'b0010001010000100001000000000000,
31'b0011000000000000000000000110000,
31'b0010001010000000001000000000000,
31'b0001000010100000000000000000000,
31'b1000000000000000010000000100010,
31'b1000000000000000000000111000000,
31'b1000000000000100010000000100010,
31'b1000000000000000100001000000100,
31'b1000000000001000010000000100010,
31'b1000000000001000000000111000000,
31'b0000000010000000010000010000100,
31'b1000000001000001000000000000001,
31'b1000000001000011000000000000001,
31'b0001010000000001000000001000000,
31'b0100000100000000100000101000000,
31'b1000000001001001000000000000001,
31'b1000010000000001000001000000010,
31'b0011000000100000000000000110000,
31'b0010100000000000010100000100000,
31'b0001000011000000000000000000000,
31'b0010000000010000000000000101000,
31'b0000001000010000000000100000000,
31'b0000001000010010000000100000000,
31'b0001000011001000000000000000000,
31'b0011000000000000001000100000000,
31'b0000001000011000000000100000000,
31'b0000000010000000000000000011000,
31'b0000001000000100000000100000000,
31'b0010000000000000000000000101000,
31'b0000001000000000000000100000000,
31'b0000001000000010000000100000000,
31'b0000000000000000101000000010000,
31'b0010000000001000000000000101000,
31'b0000001000001000000000100000000,
31'b0000001000001010000000100000000,
31'b1000000000010001000000000000001,
31'b1000000001000000010000000100010,
31'b0000001000110000000000100000000,
31'b0100000000010001000001000001000,
31'b1000000001000000100001000000100,
31'b0110000100000000000000001001000,
31'b0100001000000000000100000001010,
31'b0100000000000000000010110000000,
31'b1000000000000001000000000000001,
31'b1000000000000011000000000000001,
31'b0000001000100000000000100000000,
31'b0100000000000001000001000001000,
31'b1000000000001001000000000000001,
31'b1000010000000000100100000100000,
31'b0000001000101000000000100000000,
31'b0100000000010000000010110000000,
31'b0001000100000000000000000000000,
31'b0001000100000010000000000000000,
31'b0001000100000100000000000000000,
31'b0001000100000110000000000000000,
31'b0001000100001000000000000000000,
31'b0001000100001010000000000000000,
31'b0001000100001100000000000000000,
31'b0000100000000001000100000000000,
31'b0001000100010000000000000000000,
31'b1010000000000001000000000000010,
31'b0001000100010100000000000000000,
31'b1010000000000101000000000000010,
31'b0001000100011000000000000000000,
31'b1010000000001001000000000000010,
31'b0011000000000001000001001000000,
31'b0010001100000000001000000000000,
31'b0001000100100000000000000000000,
31'b0001000100100010000000000000000,
31'b0001000100100100000000000000000,
31'b0001000100100110000000000000000,
31'b0000000000000000000100000001100,
31'b0001100001000000000000010000000,
31'b0001000000000001010000000010000,
31'b0000100000100001000100000000000,
31'b0001000100110000000000000000000,
31'b1010000000100001000000000000010,
31'b0001010000000000000001000110000,
31'b1100000000000000000001000100010,
31'b0101000000000000000000001100000,
31'b0101000000000010000000001100000,
31'b1100000000000000110000000000100,
31'b0010001100100000001000000000000,
31'b0001000101000000000000000000000,
31'b0001000101000010000000000000000,
31'b0000100000000000010000000000100,
31'b0000100000000010010000000000100,
31'b0001000101001000000000000000000,
31'b0001100000100000000000010000000,
31'b0000100000001000010000000000100,
31'b0000000100000000000000000011000,
31'b0001000101010000000000000000000,
31'b1010000001000001000000000000010,
31'b0000100000010000010000000000100,
31'b0000111000001000000000000000001,
31'b0001000101011000000000000000000,
31'b0001100000110000000000010000000,
31'b1000010000000000000000100001100,
31'b0000111000000000000000000000001,
31'b0001000101100000000000000000000,
31'b0000000000000001010000000001000,
31'b0000100000100000010000000000100,
31'b0001000000000000000100000010100,
31'b0001100000000010000000010000000,
31'b0001100000000000000000010000000,
31'b0001100000000110000000010000000,
31'b0001100000000100000000010000000,
31'b1001000000000010000010000100000,
31'b1001000000000000000010000100000,
31'b0010101000000000001000010000000,
31'b1100000000000001100100000000000,
31'b0110110000000000000000000000100,
31'b0001100000010000000000010000000,
31'b1100010000000000000000000100001,
31'b0001100000010100000000010000000,
31'b0001000110000000000000000000000,
31'b0001000110000010000000000000000,
31'b0100100000000000000010100000000,
31'b0101000000000000100100000000001,
31'b0001000110001000000000000000000,
31'b0001110000000000000000100000001,
31'b0101010000000001000000000100000,
31'b0000100010000001000100000000000,
31'b0001000110010000000000000000000,
31'b1010000010000001000000000000010,
31'b0101000000000000010001000000000,
31'b0101000000000010010001000000000,
31'b0001010000000000010000001010000,
31'b1100000000000000010000001000010,
31'b1100000000000000000000110100000,
31'b0010001110000000001000000000000,
31'b1010000000000000000010000001000,
31'b1010000000000010000010000001000,
31'b1010000000000100000010000001000,
31'b1010010000000000000000001000010,
31'b0011010000000000000001000000000,
31'b0110000001000000000000001001000,
31'b0011010000000100000001000000000,
31'b0000101000010000000000110000000,
31'b1010000000010000000010000001000,
31'b0100000000001000000001010000100,
31'b0101000000100000010001000000000,
31'b0100000000000000100000101000000,
31'b0101000010000000000000001100000,
31'b0100000000000000000001010000100,
31'b1000000001000000100010100000000,
31'b0000101000000000000000110000000,
31'b0001000111000000000000000000000,
31'b0011000000100000000000000000011,
31'b0000100010000000010000000000100,
31'b1000100000001000000000101000000,
31'b0001010000000000001000010000010,
31'b1100000000000000001000010010000,
31'b1000100000000010000000101000000,
31'b1000100000000000000000101000000,
31'b0000000000000000010010000000010,
31'b0010000100000000000000000101000,
31'b0000001100000000000000100000000,
31'b0000010000000000010000001001000,
31'b0000000100000000101000000010000,
31'b0110000000000000001000000000110,
31'b1000000000000000010000000010001,
31'b1000100000010000000000101000000,
31'b1010000001000000000010000001000,
31'b0011000000000000000000000000011,
31'b0000100010100000010000000000100,
31'b0011000000000100000000000000011,
31'b0110000000000010000000001001000,
31'b0110000000000000000000001001000,
31'b1010000000000000000001001000001,
31'b1011000000000000000010000010000,
31'b1000000100000001000000000000001,
31'b1001000010000000000010000100000,
31'b0000001100100000000000100000000,
31'b0100000100000001000001000001000,
31'b1000000100001001000000000000001,
31'b0110000000010000000000001001000,
31'b1000000000000000100010100000000,
31'b1001100000000000000100000000001,
31'b0001001000000000000000000000000,
31'b0001001000000010000000000000000,
31'b0001001000000100000000000000000,
31'b0010000000011000001000000000000,
31'b0001001000001000000000000000000,
31'b0010000000010100001000000000000,
31'b0010000000010010001000000000000,
31'b0010000000010000001000000000000,
31'b0001001000010000000000000000000,
31'b0010000000001100001000000000000,
31'b0000000011000000000000100000000,
31'b0010000000001000001000000000000,
31'b0010000000000110001000000000000,
31'b0010000000000100001000000000000,
31'b0010000000000010001000000000000,
31'b0010000000000000001000000000000,
31'b0001001000100000000000000000000,
31'b0100010000000000011000000000000,
31'b0001001000100100000000000000000,
31'b0111000000000000000000000000101,
31'b0010010000000000000010000000100,
31'b0101000000010000000010010000000,
31'b0010010000000100000010000000100,
31'b0010000000110000001000000000000,
31'b0001001000110000000000000000000,
31'b0101000000001000000010010000000,
31'b0000010000000000000000010000001,
31'b0010000000101000001000000000000,
31'b0101000000000010000010010000000,
31'b0101000000000000000010010000000,
31'b0010000000100010001000000000000,
31'b0010000000100000001000000000000,
31'b0001001001000000000000000000000,
31'b0001001001000010000000000000000,
31'b0000000010010000000000100000000,
31'b0000001000001000000000000011000,
31'b0010000000000000000000100110000,
31'b0001000000010000100000000100000,
31'b0000001000000010000000000011000,
31'b0000001000000000000000000011000,
31'b0000000010000100000000100000000,
31'b0001000000001000100000000100000,
31'b0000000010000000000000100000000,
31'b0000000010000010000000100000000,
31'b0001000000000010100000000100000,
31'b0001000000000000100000000100000,
31'b0000000010001000000000100000000,
31'b0010000001000000001000000000000,
31'b0001001001100000000000000000000,
31'b0101000100000000100000001000000,
31'b0000001000000001000100010000000,
31'b0000001000101000000000000011000,
31'b0010010001000000000010000000100,
31'b0001101100000000000000010000000,
31'b0100000010000000000100000001010,
31'b0000001000100000000000000011000,
31'b1001000000000000000000011000000,
31'b1001000000000010000000011000000,
31'b0000000010100000000000100000000,
31'b0000000010100010000000100000000,
31'b1001000000001000000000011000000,
31'b0001000000100000100000000100000,
31'b0000000010101000000000100000000,
31'b0000000000000000000001010000010,
31'b0001001010000000000000000000000,
31'b0000000000000000001000000110000,
31'b0000000001010000000000100000000,
31'b0000000001010010000000100000000,
31'b0010000000000000100000000001000,
31'b0010000000000010100000000001000,
31'b0010000000000100100000000001000,
31'b0010000010010000001000000000000,
31'b0000000001000100000000100000000,
31'b0000000001000110000000100000000,
31'b0000000001000000000000100000000,
31'b0000000001000010000000100000000,
31'b0010000000010000100000000001000,
31'b0010000010000100001000000000000,
31'b0000000001001000000000100000000,
31'b0010000010000000001000000000000,
31'b1000010000000000000100000000000,
31'b1000010000000010000100000000000,
31'b1000010000000100000100000000000,
31'b1000010000000110000100000000000,
31'b1000010000001000000100000000000,
31'b1000010000001010000100000000000,
31'b1100100000000000100000100000000,
31'b0010100000000001100000000000100,
31'b1000010000010000000100000000000,
31'b1000010000010010000100000000000,
31'b0000000001100000000000100000000,
31'b0000010100000000001001000000000,
31'b1000010000011000000100000000000,
31'b0101000010000000000010010000000,
31'b0010110000000000000000000000010,
31'b0010000010100000001000000000000,
31'b0000000000010100000000100000000,
31'b0000000001000000001000000110000,
31'b0000000000010000000000100000000,
31'b0000000000010010000000100000000,
31'b0010000001000000100000000001000,
31'b0011001000000000001000100000000,
31'b0000000000011000000000100000000,
31'b0000001010000000000000000011000,
31'b0000000000000100000000100000000,
31'b0000000000000110000000100000000,
31'b0000000000000000000000100000000,
31'b0000000000000010000000100000000,
31'b0000000000001100000000100000000,
31'b0001000010000000100000000100000,
31'b0000000000001000000000100000000,
31'b0000000000001010000000100000000,
31'b1000010001000000000100000000000,
31'b1000010001000010000100000000000,
31'b0000000000110000000000100000000,
31'b0000000000110010000000100000000,
31'b1000010001001000000100000000000,
31'b1000010000000001010000000000100,
31'b0100000000000000000100000001010,
31'b0100001000000000000010110000000,
31'b0000000000100100000000100000000,
31'b1000000000000000000001000100100,
31'b0000000000100000000000100000000,
31'b0000000000100010000000100000000,
31'b1000000000000000110000000000010,
31'b1000000000001000000001000100100,
31'b0000000000101000000000100000000,
31'b0000000010000000000001010000010,
31'b0001001100000000000000000000000,
31'b0001001100000010000000000000000,
31'b0001001100000100000000000000000,
31'b0011000000000000000100001000010,
31'b1010000000000000000101000000000,
31'b1010000000000010000101000000000,
31'b1010000000000100000101000000000,
31'b0010000100010000001000000000000,
31'b0001001100010000000000000000000,
31'b1010001000000001000000000000010,
31'b0000100000000000000001000000010,
31'b0010000100001000001000000000000,
31'b1010000000010000000101000000000,
31'b1001100000000000000000001000000,
31'b0010000100000010001000000000000,
31'b0010000100000000001000000000000,
31'b0001001100100000000000000000000,
31'b0101000001000000100000001000000,
31'b0001001100100100000000000000000,
31'b1100010000000000100000000000001,
31'b1001000000000000100010000000000,
31'b1001000000000010100010000000000,
31'b1100000000000001000100000100000,
31'b0010000100110000001000000000000,
31'b0001100000000000100000010100000,
31'b0010000000000100000000100000011,
31'b0000100000100000000001000000010,
31'b0010000000000000000000100000011,
31'b1001000000010000100010000000000,
31'b1010000000000000000010100010000,
31'b0010010001000000000001100000000,
31'b0010000100100000001000000000000,
31'b0100000000000000010001100000000,
31'b0101000000100000100000001000000,
31'b0000101000000000010000000000100,
31'b1000010010000000000000000010100,
31'b1101000000000000000000010100000,
31'b0001101000100000000000010000000,
31'b0000110000010010000000000000001,
31'b0000110000010000000000000000001,
31'b0101100000000000000010000000000,
31'b0101100000000010000010000000000,
31'b0000000110000000000000100000000,
31'b0000110000001000000000000000001,
31'b0101100000001000000010000000000,
31'b0001000100000000100000000100000,
31'b0000110000000010000000000000001,
31'b0000110000000000000000000000001,
31'b0101000000000010100000001000000,
31'b0101000000000000100000001000000,
31'b0010100000010000001000010000000,
31'b1100000000000000010000000100100,
31'b1001000001000000100010000000000,
31'b0001101000000000000000010000000,
31'b1100000000000000100001000000010,
31'b0001101000000100000000010000000,
31'b1001000100000000000000011000000,
31'b1001001000000000000010000100000,
31'b0010100000000000001000010000000,
31'b0010100000000010001000010000000,
31'b0010010000000100000001100000000,
31'b0001101000010000000000010000000,
31'b0010010000000000000001100000000,
31'b0000110000100000000000000000001,
31'b0000000000000000000011000000100,
31'b0000000100000000001000000110000,
31'b0000000101010000000000100000000,
31'b1000010001000000000000000010100,
31'b0010000100000000100000000001000,
31'b0110000000000000011001000000000,
31'b0010000100000100100000000001000,
31'b0010000110010000001000000000000,
31'b0000000101000100000000100000000,
31'b0000010001000000000110000100000,
31'b0000000101000000000000100000000,
31'b0000010000100000001001000000000,
31'b0010000100010000100000000001000,
31'b1110000000000000000000010001000,
31'b0010000000000000000001010000001,
31'b0010000110000000001000000000000,
31'b1000010100000000000100000000000,
31'b1000010100000010000100000000000,
31'b1000010100000100000100000000000,
31'b1000000000000000000010100100000,
31'b1001000010000000100010000000000,
31'b0100000001000000010000010000010,
31'b0100100000000001000000000010010,
31'b0000100000010000000000110000000,
31'b1000010100010000000100000000000,
31'b0000010000000100001001000000000,
31'b0000010000000010001001000000000,
31'b0000010000000000001001000000000,
31'b0100000000000010001000001010000,
31'b0100000000000000001000001010000,
31'b0000100000000010000000110000000,
31'b0000100000000000000000110000000,
31'b0000000100010100000000100000000,
31'b1000010000000100000000000010100,
31'b0000000100010000000000100000000,
31'b1000010000000000000000000010100,
31'b0010000101000000100000000001000,
31'b1100000000000000000001001000100,
31'b0000000100011000000000100000000,
31'b1000101000000000000000101000000,
31'b0000000100000100000000100000000,
31'b0000010000000000000110000100000,
31'b0000000100000000000000100000000,
31'b0000000100000010000000100000000,
31'b0000000100001100000000100000000,
31'b0001100000000001000100100000000,
31'b0000000100001000000000100000000,
31'b0000110010000000000000000000001,
31'b1000010101000000000100000000000,
31'b0101000010000000100000001000000,
31'b0000000100110000000000100000000,
31'b1000010000100000000000000010100,
31'b0100000000000100000000101100000,
31'b0100000000000000010000010000010,
31'b0100000000000000000000101100000,
31'b0100000000000100010000010000010,
31'b1000000000000000001010000010000,
31'b1000000100000000000001000100100,
31'b0000000100100000000000100000000,
31'b0000010001000000001001000000000,
31'b0000000000000100001000000000011,
31'b0100000001000000001000001010000,
31'b0000000000000000001000000000011,
31'b0000100001000000000000110000000,
31'b0001010000000000000000000000000,
31'b0001010000000010000000000000000,
31'b0001010000000100000000000000000,
31'b0100000000001000000010000000001,
31'b0001010000001000000000000000000,
31'b0100000000000100000010000000001,
31'b0100000000000010000010000000001,
31'b0100000000000000000010000000001,
31'b0001010000010000000000000000000,
31'b0110000000000000000000010000100,
31'b0001010000010100000000000000000,
31'b0110000000000100000000010000100,
31'b0001010000011000000000000000000,
31'b0110000000001000000000010000100,
31'b0111000000100000010000000000000,
31'b0100000000010000000010000000001,
31'b0001010000100000000000000000000,
31'b0100001000000000011000000000000,
31'b0001010000100100000000000000000,
31'b0100001000000100011000000000000,
31'b0010001000000000000010000000100,
31'b0100001000001000011000000000000,
31'b0111000000010000010000000000000,
31'b0100000000100000000010000000001,
31'b0001010000110000000000000000000,
31'b0110000000100000000000010000100,
31'b0000001000000000000000010000001,
31'b0001000000000000001010000000100,
31'b0111000000000100010000000000000,
31'b1000000010000001000001000000010,
31'b0111000000000000010000000000000,
31'b0111000000000010010000000000000,
31'b0001010001000000000000000000000,
31'b0100000000000000000001001001000,
31'b1000000000000000000000001000001,
31'b1000000000000010000000001000001,
31'b0001010001001000000000000000000,
31'b0001000000000000000001000000011,
31'b1000000000001000000000001000001,
31'b0000010000000000000000000011000,
31'b0001010001010000000000000000000,
31'b0110000001000000000000010000100,
31'b1000000000010000000000001000001,
31'b1000100000000000010000100010000,
31'b0001010001011000000000000000000,
31'b0001011000000000100000000100000,
31'b1000000100000000000000100001100,
31'b0000101100000000000000000000001,
31'b0001010001100000000000000000000,
31'b0100001001000000011000000000000,
31'b1000000000100000000000001000001,
31'b1010000000000000100100000010000,
31'b0011100000000000000000100000010,
31'b0001110100000000000000010000000,
31'b1000000000101000000000001000001,
31'b0000010000100000000000000011000,
31'b1001000000000100000100100000000,
31'b0110000000000000010000000011000,
31'b1001000000000000000100100000000,
31'b1001000000000010000100100000000,
31'b0110100100000000000000000000100,
31'b0000100000000000100000000010010,
31'b1100000100000000000000000100001,
31'b0000101100100000000000000000001,
31'b0001010010000000000000000000000,
31'b0100100000000000000100000100000,
31'b0001010010000100000000000000000,
31'b0100100000000100000100000100000,
31'b0001010010001000000000000000000,
31'b0100100000001000000100000100000,
31'b0101000100000001000000000100000,
31'b0100000010000000000010000000001,
31'b0001010010010000000000000000000,
31'b0110000010000000000000010000100,
31'b0001000000100001000000001000000,
31'b0001010000000000101000000001000,
31'b0001010010011000000000000000000,
31'b1100000000000000000110010000000,
31'b0011010000000000000000000110000,
31'b1110000000000000000000000100010,
31'b1000001000000000000100000000000,
31'b1000001000000010000100000000000,
31'b1000001000000100000100000000000,
31'b1010000100000000000000001000010,
31'b1000001000001000000100000000000,
31'b1000001000001010000100000000000,
31'b1000100000000000001001001000000,
31'b0100000010100000000010000000001,
31'b1000001000010000000100000000000,
31'b1000001000010010000100000000000,
31'b0001000000000001000000001000000,
31'b0001000000000011000000001000000,
31'b1000001000011000000100000000000,
31'b1000000000000001000001000000010,
31'b0010101000000000000000000000010,
31'b1011000000000000001100000000000,
31'b0001010011000000000000000000000,
31'b0100100001000000000100000100000,
31'b1000000010000000000000001000001,
31'b1000001100000000000000000010100,
31'b0001010011001000000000000000000,
31'b0011010000000000001000100000000,
31'b1000101000000000010000000001000,
31'b0000010010000000000000000011000,
31'b0000000000000000000100011000000,
31'b0010010000000000000000000101000,
31'b0000011000000000000000100000000,
31'b0000011000000010000000100000000,
31'b0000010000000000101000000010000,
31'b1010000000000001001000010000000,
31'b0000100000000000000000001010100,
31'b0000101110000000000000000000001,
31'b1000001001000000000100000000000,
31'b1000001001000010000100000000000,
31'b1000001001000100000100000000000,
31'b0100100000000000001011000000000,
31'b1000001001001000000100000000000,
31'b1000001000000001010000000000100,
31'b0110000100000000000010000000010,
31'b0100000000000000010000000101000,
31'b1000010000000001000000000000001,
31'b1000010000000011000000000000001,
31'b0001000001000001000000001000000,
31'b0101000000000000011000100000000,
31'b1000010000001001000000000000001,
31'b1000000000000000100100000100000,
31'b0011000000000000000010100000100,
31'b1101000000000001000010000000000,
31'b0001010100000000000000000000000,
31'b0100000000000001100000100000000,
31'b0001010100000100000000000000000,
31'b0100000100001000000010000000001,
31'b0001010100001000000000000000000,
31'b0100000100000100000010000000001,
31'b0101000010000001000000000100000,
31'b0100000100000000000010000000001,
31'b0001010100010000000000000000000,
31'b1010010000000001000000000000010,
31'b0001010100010100000000000000000,
31'b0000101001001000000000000000001,
31'b0001010100011000000000000000000,
31'b0000101001000100000000000000001,
31'b1000000001000000000000100001100,
31'b0000101001000000000000000000001,
31'b0001010100100000000000000000000,
31'b0100001100000000011000000000000,
31'b0001010100100100000000000000000,
31'b1100001000000000100000000000001,
31'b0011000010000000000001000000000,
31'b0011000010000010000001000000000,
31'b0011000010000100000001000000000,
31'b1100000000000001010000000000010,
31'b0001010100110000000000000000000,
31'b0000100010001000000100001000000,
31'b0001000000000000000001000110000,
31'b0000001010000000001001000000000,
31'b0110100001000000000000000000100,
31'b0000100010000000000100001000000,
31'b1100000001000000000000000100001,
31'b0000101001100000000000000000001,
31'b0001010101000000000000000000000,
31'b0100000100000000000001001001000,
31'b1000000100000000000000001000001,
31'b1000001010000000000000000010100,
31'b0001010101001000000000000000000,
31'b0001110000100000000000010000000,
31'b1000000100001000000000001000001,
31'b0000101000010000000000000000001,
31'b0001010101010000000000000000000,
31'b0000101000001100000000000000001,
31'b1000000100010000000000001000001,
31'b0000101000001000000000000000001,
31'b1010000000000001000001000000001,
31'b0000101000000100000000000000001,
31'b1000000000000000000000100001100,
31'b0000101000000000000000000000001,
31'b0001010101100000000000000000000,
31'b0001000000000000001001100000000,
31'b1100000000000000000100000000110,
31'b0010000010000000000001000011000,
31'b0110100000010000000000000000100,
31'b0001110000000000000000010000000,
31'b1100000000010000000000000100001,
31'b0001110000000100000000010000000,
31'b0110100000001000000000000000100,
31'b0000100000000000011010000000000,
31'b1100000000001000000000000100001,
31'b0000101000101000000000000000001,
31'b0110100000000000000000000000100,
31'b0000000000000000000001000101000,
31'b1100000000000000000000000100001,
31'b0000101000100000000000000000001,
31'b0001010110000000000000000000000,
31'b0100100100000000000100000100000,
31'b0101000000001001000000000100000,
31'b1010000000100000000000001000010,
31'b0000000000000000100110000000000,
31'b0001100000000000000000100000001,
31'b0101000000000001000000000100000,
31'b0101000000000011000000000100000,
31'b0001010110010000000000000000000,
31'b0000100000101000000100001000000,
31'b0101010000000000010001000000000,
31'b0000001000100000001001000000000,
31'b0001000000000000010000001010000,
31'b0000100000100000000100001000000,
31'b1100000000000000010010000001000,
31'b0000101011000000000000000000001,
31'b1000001100000000000100000000000,
31'b1010000000000100000000001000010,
31'b1010000000000010000000001000010,
31'b1010000000000000000000001000010,
31'b0011000000000000000001000000000,
31'b0011000000000010000001000000000,
31'b0011000000000100000001000000000,
31'b1010000000001000000000001000010,
31'b1010100000000001001000000000000,
31'b0000100000001000000100001000000,
31'b0001000100000001000000001000000,
31'b0000001000000000001001000000000,
31'b0011000000010000000001000000000,
31'b0000100000000000000100001000000,
31'b0011000000010100000001000000000,
31'b0000100000000100000100001000000,
31'b0001010111000000000000000000000,
31'b1100000000000000100100001000000,
31'b1000001000000010000000000010100,
31'b1000001000000000000000000010100,
31'b0001000000000000001000010000010,
31'b1000101000000000000100010000000,
31'b0110000000100000000010000000010,
31'b1000110000000000000000101000000,
31'b0000010000000000010010000000010,
31'b0000001000000000000110000100000,
31'b0000011100000000000000100000000,
31'b0000000000000000010000001001000,
31'b0001000001000000010000001010000,
31'b0000101010000100000000000000001,
31'b1000010000000000010000000010001,
31'b0000101010000000000000000000001,
31'b1110000000000000000000000010001,
31'b0011010000000000000000000000011,
31'b0110000000001000000010000000010,
31'b0010000000000000000001000011000,
31'b0100000000000000000100010100000,
31'b0110010000000000000000001001000,
31'b0110000000000000000010000000010,
31'b0110000000000010000010000000010,
31'b1100100000000000000110000000000,
31'b0000100010000000011010000000000,
31'b0001000101000001000000001000000,
31'b0000001001000000001001000000000,
31'b0110100010000000000000000000100,
31'b0000100001000000000100001000000,
31'b1100000010000000000000000100001,
31'b0000101010100000000000000000001,
31'b0001011000000000000000000000000,
31'b0100000000100000011000000000000,
31'b0001011000000100000000000000000,
31'b0100001000001000000010000000001,
31'b0010000000100000000010000000100,
31'b0100001000000100000010000000001,
31'b0101000000000000001000010000100,
31'b0100001000000000000010000000001,
31'b0001011000010000000000000000000,
31'b0110001000000000000000010000100,
31'b0000000000100000000000010000001,
31'b0010010000001000001000000000000,
31'b0010010000000110001000000000000,
31'b0010010000000100001000000000000,
31'b0010010000000010001000000000000,
31'b0010010000000000001000000000000,
31'b1000000010000000000100000000000,
31'b0100000000000000011000000000000,
31'b0000000000010000000000010000001,
31'b0100000000000100011000000000000,
31'b0010000000000000000010000000100,
31'b0100000000001000011000000000000,
31'b0010000000000100000010000000100,
31'b0100001000100000000010000000001,
31'b0000000000000100000000010000001,
31'b0100000000010000011000000000000,
31'b0000000000000000000000010000001,
31'b0000000000000010000000010000001,
31'b0010000000010000000010000000100,
31'b0101010000000000000010010000000,
31'b0000000000001000000000010000001,
31'b0010010000100000001000000000000,
31'b0001011001000000000000000000000,
31'b0100001000000000000001001001000,
31'b1000001000000000000000001000001,
31'b1000001000000010000000001000001,
31'b0010010000000000000000100110000,
31'b0001010000010000100000000100000,
31'b1000100010000000010000000001000,
31'b0000100100010000000000000000001,
31'b0001000000000001000100000000001,
31'b0001010000001000100000000100000,
31'b0000010010000000000000100000000,
31'b0000100100001000000000000000001,
31'b0100100010000000100100000000000,
31'b0001010000000000100000000100000,
31'b0000100100000010000000000000001,
31'b0000100100000000000000000000001,
31'b0000000000000001000000101000000,
31'b0100000001000000011000000000000,
31'b0000000001010000000000010000001,
31'b0100100000000000000000001100001,
31'b0010000001000000000010000000100,
31'b1010000000000000001100100000000,
31'b0010000100010000000001100000000,
31'b0001100000000000000000000101010,
31'b0000000001000100000000010000001,
31'b0100000001010000011000000000000,
31'b0000000001000000000000010000001,
31'b0000100000000000001000100000010,
31'b0010000100000100000001100000000,
31'b0001010000100000100000000100000,
31'b0010000100000000000001100000000,
31'b0000100100100000000000000000001,
31'b1000000000100000000100000000000,
31'b1000000000100010000100000000000,
31'b1000000000100100000100000000000,
31'b1000000101000000000000000010100,
31'b1000000000101000000100000000000,
31'b1000000000101010000100000000000,
31'b1000100001000000010000000001000,
31'b0100001010000000000010000000001,
31'b1000000000110000000100000000000,
31'b1000000000110010000100000000000,
31'b0000010001000000000000100000000,
31'b0000010001000010000000100000000,
31'b1100000000000000000000100001010,
31'b0010010010000100001000000000000,
31'b0010100000100000000000000000010,
31'b0010010010000000001000000000000,
31'b1000000000000000000100000000000,
31'b1000000000000010000100000000000,
31'b1000000000000100000100000000000,
31'b1000000000000110000100000000000,
31'b1000000000001000000100000000000,
31'b1000000000001010000100000000000,
31'b1000000000001100000100000000000,
31'b1001100100000001000000000000000,
31'b1000000000010000000100000000000,
31'b1000000000010010000100000000000,
31'b0000000010000000000000010000001,
31'b0000000100000000001001000000000,
31'b1000000000011000000100000000000,
31'b1000001000000001000001000000010,
31'b0010100000000000000000000000010,
31'b0010100000000010000000000000010,
31'b1000000001100000000100000000000,
31'b1000000100000100000000000010100,
31'b0000010000010000000000100000000,
31'b1000000100000000000000000010100,
31'b1000100000000100010000000001000,
31'b1000100100000000000100010000000,
31'b1000100000000000010000000001000,
31'b1000100000000010010000000001000,
31'b0000010000000100000000100000000,
31'b0000010000000110000000100000000,
31'b0000010000000000000000100000000,
31'b0000010000000010000000100000000,
31'b0100100000000000100100000000000,
31'b0101000000000000000010100000001,
31'b0000010000001000000000100000000,
31'b0000100110000000000000000000001,
31'b1000000001000000000100000000000,
31'b1000000001000010000100000000000,
31'b1000000001000100000100000000000,
31'b1000000100100000000000000010100,
31'b1000000001001000000100000000000,
31'b1000000000000001010000000000100,
31'b1000100000100000010000000001000,
31'b1001000000000000000100000011000,
31'b1000000001010000000100000000000,
31'b1000010000000000000001000100100,
31'b0000010000100000000000100000000,
31'b0000010000100010000000100000000,
31'b1000010000000000110000000000010,
31'b1000001000000000100100000100000,
31'b0010100001000000000000000000010,
31'b0010100001000010000000000000010,
31'b0001011100000000000000000000000,
31'b0100001000000001100000100000000,
31'b0001011100000100000000000000000,
31'b1100000000100000100000000000001,
31'b1010010000000000000101000000000,
31'b0100000000000101001000000010000,
31'b0100000000000011001000000010000,
31'b0100000000000001001000000010000,
31'b0001100000000000000000000011001,
31'b0000100001001100000000000000001,
31'b0000110000000000000001000000010,
31'b0000100001001000000000000000001,
31'b0100100000000000000000001010010,
31'b0000100001000100000000000000001,
31'b0000100001000010000000000000001,
31'b0000100001000000000000000000001,
31'b0000000000000000100001000001000,
31'b0100000100000000011000000000000,
31'b0000000100010000000000010000001,
31'b1100000000000000100000000000001,
31'b0010000100000000000010000000100,
31'b0100000100001000011000000000000,
31'b0010000100000100000010000000100,
31'b1100000000001000100000000000001,
31'b0000000100000100000000010000001,
31'b0000000010000100001001000000000,
31'b0000000100000000000000010000001,
31'b0000000010000000001001000000000,
31'b0010000100010000000010000000100,
31'b0000101010000000000100001000000,
31'b0010000001000000000001100000000,
31'b0000100001100000000000000000001,
31'b0101000000000001001000000001000,
31'b1010000000000000000100000000011,
31'b1000001100000000000000001000001,
31'b1000000010000000000000000010100,
31'b0100100000000000011000010000000,
31'b0000100000010100000000000000001,
31'b0000100000010010000000000000001,
31'b0000100000010000000000000000001,
31'b0101110000000000000010000000000,
31'b0000100000001100000000000000001,
31'b0000100000001010000000000000001,
31'b0000100000001000000000000000001,
31'b0100000000000001000000100100000,
31'b0000100000000100000000000000001,
31'b0000100000000010000000000000001,
31'b0000100000000000000000000000001,
31'b0000000100000001000000101000000,
31'b0101010000000000100000001000000,
31'b0010000000011000000001100000000,
31'b1100000001000000100000000000001,
31'b0010000101000000000010000000100,
31'b0001111000000000000000010000000,
31'b0010000000010000000001100000000,
31'b0001000000000000100001000010000,
31'b0010000000001100000001100000000,
31'b0000101000000000011010000000000,
31'b0010000000001000000001100000000,
31'b0000100000101000000000000000001,
31'b0010000000000100000001100000000,
31'b0000100000100100000000000000001,
31'b0010000000000000000001100000000,
31'b0000100000100000000000000000001,
31'b1000000100100000000100000000000,
31'b1000000100100010000100000000000,
31'b1000000100100100000100000000000,
31'b1000000001000000000000000010100,
31'b1001000000000000000000000001100,
31'b1001000000000010000000000001100,
31'b1001000000000100000000000001100,
31'b1001100000100001000000000000000,
31'b1000000100110000000100000000000,
31'b0000000001000000000110000100000,
31'b0000010101000000000000100000000,
31'b0000000000100000001001000000000,
31'b1100000000000000000100001100000,
31'b0000101000100000000100001000000,
31'b0010100100100000000000000000010,
31'b0000100011000000000000000000001,
31'b1000000100000000000100000000000,
31'b1000000100000010000100000000000,
31'b1000000100000100000100000000000,
31'b0000000000010000001001000000000,
31'b1000000100001000000100000000000,
31'b1001100000000101000000000000000,
31'b1001100000000011000000000000000,
31'b1001100000000001000000000000000,
31'b1000000100010000000100000000000,
31'b0000000000000100001001000000000,
31'b0000000000000010001001000000000,
31'b0000000000000000001001000000000,
31'b1001000000000000001000001000010,
31'b0000101000000000000100001000000,
31'b0010100100000000000000000000010,
31'b0000000000001000001001000000000,
31'b1000000101100000000100000000000,
31'b1000000000000100000000000010100,
31'b1000000000000010000000000010100,
31'b1000000000000000000000000010100,
31'b1001000001000000000000000001100,
31'b1000100000000000000100010000000,
31'b1000100100000000010000000001000,
31'b1000000000001000000000000010100,
31'b0000010100000100000000100000000,
31'b0000000000000000000110000100000,
31'b0000010100000000000000100000000,
31'b0010000000000000000000010000010,
31'b0100100100000000100100000000000,
31'b0000100010000100000000000000001,
31'b0000100010000010000000000000001,
31'b0000100010000000000000000000001,
31'b1000000101000000000100000000000,
31'b1000000101000010000100000000000,
31'b1000000101000100000100000000000,
31'b1000000000100000000000000010100,
31'b1001000000000000010000010010000,
31'b1000100000100000000100010000000,
31'b0110001000000000000010000000010,
31'b1001100001000001000000000000000,
31'b1000010000000000001010000010000,
31'b0000000001000100001001000000000,
31'b0000010100100000000000100000000,
31'b0000000001000000001001000000000,
31'b0011000000000000010000000000110,
31'b0000101001000000000100001000000,
31'b0010000010000000000001100000000,
31'b0000100010100000000000000000001,
31'b0001100000000000000000000000000,
31'b0001100000000010000000000000000,
31'b0001100000000100000000000000000,
31'b0001100000000110000000000000000,
31'b0001100000001000000000000000000,
31'b0001100000001010000000000000000,
31'b0001100000001100000000000000000,
31'b0000000100000001000100000000000,
31'b0001100000010000000000000000000,
31'b0010000000000000000101001000000,
31'b0001100000010100000000000000000,
31'b0010101000001000001000000000000,
31'b1000000000000001001001000000000,
31'b1001001100000000000000001000000,
31'b1011000000000000000100000000010,
31'b0010101000000000001000000000000,
31'b0001100000100000000000000000000,
31'b0000000000000000010100000010000,
31'b0001100000100100000000000000000,
31'b0001000000000001000000000001100,
31'b0001100000101000000000000000000,
31'b0001000101000000000000010000000,
31'b0001100000101100000000000000000,
31'b0000100000000000010000010000100,
31'b0001100000110000000000000000000,
31'b0001000000000000100010001000000,
31'b0001100000110100000000000000000,
31'b1100000000000000100000000011000,
31'b1101000001000000100000000000000,
31'b0001000101010000000000010000000,
31'b1110000000000000001000000100000,
31'b0010101000100000001000000000000,
31'b0001100001000000000000000000000,
31'b0001100001000010000000000000000,
31'b0000000100000000010000000000100,
31'b0000100000001000000000000011000,
31'b0001100001001000000000000000000,
31'b0001000100100000000000010000000,
31'b0000100000000010000000000011000,
31'b0000100000000000000000000011000,
31'b0100000010000000000001000000100,
31'b0101000000000000000000011100000,
31'b0000101010000000000000100000000,
31'b1000010000000000010000100010000,
31'b1101000000100000100000000000000,
31'b0001101000000000100000000100000,
31'b0000101010001000000000100000000,
31'b0000100000010000000000000011000,
31'b0001100001100000000000000000000,
31'b0001000100001000000000010000000,
31'b0000100000000001000100010000000,
31'b0001000100001100000000010000000,
31'b0000000000000001000000000010100,
31'b0001000100000000000000010000000,
31'b0001000000000000010100000001000,
31'b0001000100000100000000010000000,
31'b1101000000001000100000000000000,
31'b0001000100011000000000010000000,
31'b0010001100000000001000010000000,
31'b1100000010000000000000100100000,
31'b1101000000000000100000000000000,
31'b0001000100010000000000010000000,
31'b1101000000000100100000000000000,
31'b0001000100010100000000010000000,
31'b0001100010000000000000000000000,
31'b0100010000000000000100000100000,
31'b0100000100000000000010100000000,
31'b0100010000000100000100000100000,
31'b0100000000000001100000000000001,
31'b0100010000001000000100000100000,
31'b0100000100001000000010100000000,
31'b0000100000000000100000100100000,
31'b0100000001000000000001000000100,
31'b0100010000010000000100000100000,
31'b0001000000000000000010000000110,
31'b1000000001000000000000000001101,
31'b1001000000000000000000000010101,
31'b1000000100000001000000010000001,
31'b0011100000000000000000000110000,
31'b0010101010000000001000000000000,
31'b1100000000000000001000000010000,
31'b0001010000000000001000000000010,
31'b1100000000000100001000000010000,
31'b0010010000000001000101000000000,
31'b1100000000001000001000000010000,
31'b0001010000001000001000000000010,
31'b1100001000000000100000100000000,
31'b0010001000000001100000000000100,
31'b1100000000010000001000000010000,
31'b0001010000010000001000000000010,
31'b0010011000001000000000000000010,
31'b1100000001000000000000100100000,
31'b0010011000000100000000000000010,
31'b0000010100000000000100001000000,
31'b0010011000000000000000000000010,
31'b0010000000000000010100000100000,
31'b0100000000010000000001000000100,
31'b0100010001000000000100000100000,
31'b0000101000010000000000100000000,
31'b1000000100001000000000101000000,
31'b0100000001000001100000000000001,
31'b1010000000000000000010010001000,
31'b1000011000000000010000000001000,
31'b1000000100000000000000101000000,
31'b0100000000000000000001000000100,
31'b0100000000000010000001000000100,
31'b0000101000000000000000100000000,
31'b1000000000000000000000000001101,
31'b0100000000001000000001000000100,
31'b0100000000001010000001000000100,
31'b0000101000001000000000100000000,
31'b1000000100010000000000101000000,
31'b1100000001000000001000000010000,
31'b0001010001000000001000000000010,
31'b0010001000000000110100000000000,
31'b1100000000010000000000100100000,
31'b0001000000000000001001000000001,
31'b0001000110000000000000010000000,
31'b0010010000000000010001000000100,
31'b1101000000000000001000000001000,
31'b1000100000000001000000000000001,
31'b1100000000000100000000100100000,
31'b0010000000000001000000000100100,
31'b1100000000000000000000100100000,
31'b1101000010000000100000000000000,
31'b0001000110010000000000010000000,
31'b0010011001000000000000000000010,
31'b1100000000001000000000100100000,
31'b0001100100000000000000000000000,
31'b0001100100000010000000000000000,
31'b0000000001000000010000000000100,
31'b0000000000001001000100000000000,
31'b0001100100001000000000000000000,
31'b0000000000000101000100000000000,
31'b0000000000000011000100000000000,
31'b0000000000000001000100000000000,
31'b0001100100010000000000000000000,
31'b1010100000000001000000000000010,
31'b0000001000000000000001000000010,
31'b0000001000000010000001000000010,
31'b1001001000000010000000001000000,
31'b1001001000000000000000001000000,
31'b0000001000001000000001000000010,
31'b0000000000010001000100000000000,
31'b0001100100100000000000000000000,
31'b0001000001001000000000010000000,
31'b0000000000000000000000010011000,
31'b0000000000101001000100000000000,
31'b0001000001000010000000010000000,
31'b0001000001000000000000010000000,
31'b0000000000100011000100000000000,
31'b0000000000100001000100000000000,
31'b0001100100110000000000000000000,
31'b0001000100000000100010001000000,
31'b0000001000100000000001000000010,
31'b0100000010000000000101000010000,
31'b0110010001000000000000000000100,
31'b0001000001010000000000010000000,
31'b0000001010000010000000110000000,
31'b0000001010000000000000110000000,
31'b0000000000000100010000000000100,
31'b0001000000101000000000010000000,
31'b0000000000000000010000000000100,
31'b0000000000000010010000000000100,
31'b0001000000100010000000010000000,
31'b0001000000100000000000010000000,
31'b0000000000001000010000000000100,
31'b0000000001000001000100000000000,
31'b0101001000000000000010000000000,
31'b0101001000000010000010000000000,
31'b0000000000010000010000000000100,
31'b0000011000001000000000000000001,
31'b0110010000100000000000000000100,
31'b0001000000110000000000010000000,
31'b0000011000000010000000000000001,
31'b0000011000000000000000000000001,
31'b0001000000001010000000010000000,
31'b0001000000001000000000010000000,
31'b0000000000100000010000000000100,
31'b0001000000001100000000010000000,
31'b0001000000000010000000010000000,
31'b0001000000000000000000010000000,
31'b0001000000000110000000010000000,
31'b0001000000000100000000010000000,
31'b0110010000001000000000000000100,
31'b0001000000011000000000010000000,
31'b0010001000000000001000010000000,
31'b0011000000000000000010000000101,
31'b0110010000000000000000000000100,
31'b0001000000010000000000010000000,
31'b0110010000000100000000000000100,
31'b0001000000010100000000010000000,
31'b0100000000000100000010100000000,
31'b0100010100000000000100000100000,
31'b0100000000000000000010100000000,
31'b0100000000000010000010100000000,
31'b0100000100000001100000000000001,
31'b0001010000000000000000100000001,
31'b0100000000001000000010100000000,
31'b0000000010000001000100000000000,
31'b0100000101000000000001000000100,
31'b1010000000000000100000001001000,
31'b0100000000010000000010100000000,
31'b0100000000100000000101000010000,
31'b1000000000000011000000010000001,
31'b1000000000000001000000010000001,
31'b0100000000011000000010100000000,
31'b0000001000100000000000110000000,
31'b1100000100000000001000000010000,
31'b0001010100000000001000000000010,
31'b0100000000100000000010100000000,
31'b0100000000100010000010100000000,
31'b0011110000000000000001000000000,
31'b0001000011000000000000010000000,
31'b0100001000000001000000000010010,
31'b0000001000010000000000110000000,
31'b1010010000000001001000000000000,
31'b0000010000001000000100001000000,
31'b0100000000110000000010100000000,
31'b0100000000000000000101000010000,
31'b0010000000000000000000010101000,
31'b0000010000000000000100001000000,
31'b0000001000000010000000110000000,
31'b0000001000000000000000110000000,
31'b0001000000000000000001100000010,
31'b1000000000001100000000101000000,
31'b0000000010000000010000000000100,
31'b1000000000001000000000101000000,
31'b1000000000000110000000101000000,
31'b1000000000000100000000101000000,
31'b1000000000000010000000101000000,
31'b1000000000000000000000101000000,
31'b0100000100000000000001000000100,
31'b0100000100000010000001000000100,
31'b0000101100000000000000100000000,
31'b1000000100000000000000000001101,
31'b0110000000000000100010000001000,
31'b1000000001000001000000010000001,
31'b1000100000000000010000000010001,
31'b1000000000010000000000101000000,
31'b0001000010001010000000010000000,
31'b0001000010001000000000010000000,
31'b0000000010100000010000000000100,
31'b1001000000000000000000000100110,
31'b0001000010000010000000010000000,
31'b0001000010000000000000010000000,
31'b1001000000000000110001000000000,
31'b1000000000100000000000101000000,
31'b1100010000000000000110000000000,
31'b0001000010011000000000010000000,
31'b0010001010000000001000010000000,
31'b1100000100000000000000100100000,
31'b0110010010000000000000000000100,
31'b0001000010010000000000010000000,
31'b1001000000000010000100000000001,
31'b1001000000000000000100000000001,
31'b0001101000000000000000000000000,
31'b1000000000000000001100000000010,
31'b0001101000000100000000000000000,
31'b1011000000000001000001000000000,
31'b0010000000000001000000001000010,
31'b1001000100010000000000001000000,
31'b0010100000010010001000000000000,
31'b0010100000010000001000000000000,
31'b0001101000010000000000000000000,
31'b1001000100001000000000001000000,
31'b0000000100000000000001000000010,
31'b0010100000001000001000000000000,
31'b1001000100000010000000001000000,
31'b1001000100000000000000001000000,
31'b0010100000000010001000000000000,
31'b0010100000000000001000000000000,
31'b0001101000100000000000000000000,
31'b1101000000000000000000000100000,
31'b0001101000100100000000000000000,
31'b1101000000000100000000000100000,
31'b0010110000000000000010000000100,
31'b1101000000001000000000000100000,
31'b1100000010000000100000100000000,
31'b0010100000110000001000000000000,
31'b0001101000110000000000000000000,
31'b1101000000010000000000000100000,
31'b0000110000000000000000010000001,
31'b0010100000101000001000000000000,
31'b0010010010000100000000000000010,
31'b1100000000000000001000100001000,
31'b0010010010000000000000000000010,
31'b0010100000100000001000000000000,
31'b0001101001000000000000000000000,
31'b1001000000000000100010010000000,
31'b0000100010010000000000100000000,
31'b0000101000001000000000000011000,
31'b0010100000000000000000100110000,
31'b0001100000010000100000000100000,
31'b1000010010000000010000000001000,
31'b0000101000000000000000000011000,
31'b0101000100000000000010000000000,
31'b0101000100000010000010000000000,
31'b0000100010000000000000100000000,
31'b0000100010000010000000100000000,
31'b0101000100001000000010000000000,
31'b0001100000000000100000000100000,
31'b0000100010001000000000100000000,
31'b0000010100000000000000000000001,
31'b0001101001100000000000000000000,
31'b1101000001000000000000000100000,
31'b0010000100010000001000010000000,
31'b1110000000000000101000000000000,
31'b0001000000000000000010001100000,
31'b0001001100000000000000010000000,
31'b1100000000000000000000000111000,
31'b0001010000000000000000000101010,
31'b1110000010000000000000000001000,
31'b0010000010000100000001000000001,
31'b0010000100000000001000010000000,
31'b0010000010000000000001000000001,
31'b1101001000000000100000000000000,
31'b0001100000100000100000000100000,
31'b0010010011000000000000000000010,
31'b0000100000000000000001010000010,
31'b0100000000000000010000000000010,
31'b0100000000000010010000000000010,
31'b0100000000000100010000000000010,
31'b0100000000000110010000000000010,
31'b0100000000001000010000000000010,
31'b0100000000001010010000000000010,
31'b1100000000100000100000100000000,
31'b0010100010010000001000000000000,
31'b0100000000010000010000000000010,
31'b0100000001000001000000000100001,
31'b0000100001000000000000100000000,
31'b0000100001000010000000100000000,
31'b0100010001000000100100000000000,
31'b1001000110000000000000001000000,
31'b0010010000100000000000000000010,
31'b0010100010000000001000000000000,
31'b1000110000000000000100000000000,
31'b1101000010000000000000000100000,
31'b1100000000001000100000100000000,
31'b0010000001010000000001000000001,
31'b1100000000000100100000100000000,
31'b0010000000010000000010001001000,
31'b1100000000000000100000100000000,
31'b0010000000000001100000000000100,
31'b1110000001000000000000000001000,
31'b0010000001000100000001000000001,
31'b0010010000001000000000000000010,
31'b0010000001000000000001000000001,
31'b0010010000000100000000000000010,
31'b0010000000000000000010001001000,
31'b0010010000000000000000000000010,
31'b0000000100000000000000110000000,
31'b0100000001000000010000000000010,
31'b0100000001000010010000000000010,
31'b0000100000010000000000100000000,
31'b0000100000010010000000100000000,
31'b1010000000000000000100100000010,
31'b1000010100000000000100010000000,
31'b1000010000000000010000000001000,
31'b1000010000000010010000000001000,
31'b0000100000000100000000100000000,
31'b0100000000000001000000000100001,
31'b0000100000000000000000100000000,
31'b0000100000000010000000100000000,
31'b0100010000000000100100000000000,
31'b0100010000000010100100000000000,
31'b0000100000001000000000100000000,
31'b0000100000001010000000100000000,
31'b1110000000010000000000000001000,
31'b0010000100000000100000010001000,
31'b0010000000000000110100000000000,
31'b0010000000010000000001000000001,
31'b0001001000000000001001000000001,
31'b0000000100000001000000001000001,
31'b1100000001000000100000100000000,
31'b0010000001000001100000000000100,
31'b1110000000000000000000000001000,
31'b0010000000000100000001000000001,
31'b0000100000100000000000100000000,
31'b0010000000000000000001000000001,
31'b1110000000001000000000000001000,
31'b0010000001000000000010001001000,
31'b0010010001000000000000000000010,
31'b0010000000001000000001000000001,
31'b0001101100000000000000000000000,
31'b1001000000011000000000001000000,
31'b0000000000010000000001000000010,
31'b0000001000001001000100000000000,
31'b1010100000000000000101000000000,
31'b1001000000010000000000001000000,
31'b0000001000000011000100000000000,
31'b0000001000000001000100000000000,
31'b0000000000000100000001000000010,
31'b1001000000001000000000001000000,
31'b0000000000000000000001000000010,
31'b0000000000000010000001000000010,
31'b1001000000000010000000001000000,
31'b1001000000000000000000001000000,
31'b0000000000001000000001000000010,
31'b0000010001000000000000000000001,
31'b0001101100100000000000000000000,
31'b1101000100000000000000000100000,
31'b0000001000000000000000010011000,
31'b0000001000101001000100000000000,
31'b1001100000000000100010000000000,
31'b1000000000000000000100100000001,
31'b0100000010000001000000000010010,
31'b0000001000100001000100000000000,
31'b0001000000000000100000010100000,
31'b1001000000101000000000001000000,
31'b0000000000100000000001000000010,
31'b0000000010001000000000110000000,
31'b1001000000100010000000001000000,
31'b1001000000100000000000001000000,
31'b0000000010000010000000110000000,
31'b0000000010000000000000110000000,
31'b0101000000010000000010000000000,
31'b0110000000100000010000000000001,
31'b0000001000000000010000000000100,
31'b0000010000011000000000000000001,
31'b0101000000011000000010000000000,
31'b0001001000100000000000010000000,
31'b0000010000010010000000000000001,
31'b0000010000010000000000000000001,
31'b0101000000000000000010000000000,
31'b0101000000000010000010000000000,
31'b0000000001000000000001000000010,
31'b0000010000001000000000000000001,
31'b0101000000001000000010000000000,
31'b0000010000000100000000000000001,
31'b0000010000000010000000000000001,
31'b0000010000000000000000000000001,
31'b0110000000000010010000000000001,
31'b0110000000000000010000000000001,
31'b0010000000010000001000010000000,
31'b0110000000000100010000000000001,
31'b0001001000000010000000010000000,
31'b0001001000000000000000010000000,
31'b0011010000000000010010000000000,
31'b0001001000000100000000010000000,
31'b0101000000100000000010000000000,
31'b0110000000010000010000000000001,
31'b0010000000000000001000010000000,
31'b0010000000000010001000010000000,
31'b0110011000000000000000000000100,
31'b0001001000010000000000010000000,
31'b0010000000001000001000010000000,
31'b0000010000100000000000000000001,
31'b0100000100000000010000000000010,
31'b0110000000000000000010000101000,
31'b0100001000000000000010100000000,
31'b0100001000000010000010100000000,
31'b0100000100001000010000000000010,
31'b1001000010010000000000001000000,
31'b0100001000001000000010100000000,
31'b0000001010000001000100000000000,
31'b0001000000000000010000100000100,
31'b1001000010001000000000001000000,
31'b0000000010000000000001000000010,
31'b0000000010000010000001000000010,
31'b1001000010000010000000001000000,
31'b1001000010000000000000001000000,
31'b0000000010001000000001000000010,
31'b0000000000100000000000110000000,
31'b1100000000000001000010000000001,
31'b0010000001000000100000010001000,
31'b0100001000100000000010100000000,
31'b0000000000011000000000110000000,
31'b0100000000000101000000000010010,
31'b0000000001000001000000001000001,
31'b0100000000000001000000000010010,
31'b0000000000010000000000110000000,
31'b0001000010000000100000010100000,
31'b0000000000001100000000110000000,
31'b0000000010100000000001000000010,
31'b0000000000001000000000110000000,
31'b0000000000000110000000110000000,
31'b0000000000000100000000110000000,
31'b0000000000000010000000110000000,
31'b0000000000000000000000110000000,
31'b0101000010010000000010000000000,
31'b1000010000001000000100010000000,
31'b0000100100010000000000100000000,
31'b1000110000000000000000000010100,
31'b1010000000000000000000001101000,
31'b1000010000000000000100010000000,
31'b1000010100000000010000000001000,
31'b1000001000000000000000101000000,
31'b0101000010000000000010000000000,
31'b0101000010000010000010000000000,
31'b0000100100000000000000100000000,
31'b0000100100000010000000100000000,
31'b0101000010001000000010000000000,
31'b0001000000000001000100100000000,
31'b0000100100001000000000100000000,
31'b0000010010000000000000000000001,
31'b1010000000000000001100000000001,
31'b0010000000000000100000010001000,
31'b0010000100000000110100000000000,
31'b0010000100010000000001000000001,
31'b0000000000000011000000001000001,
31'b0000000000000001000000001000001,
31'b0100100000000000000000101100000,
31'b0000000001010000000000110000000,
31'b1110000100000000000000000001000,
31'b0010000100000100000001000000001,
31'b0010000010000000001000010000000,
31'b0010000100000000000001000000001,
31'b0000100000000100001000000000011,
31'b0000000001000100000000110000000,
31'b0000100000000000001000000000011,
31'b0000000001000000000000110000000,
31'b0001110000000000000000000000000,
31'b0100000010000000000100000100000,
31'b0001110000000100000000000000000,
31'b0100100000001000000010000000001,
31'b0001110000001000000000000000000,
31'b0100100000000100000010000000001,
31'b0101000000000000100100100000000,
31'b0100100000000000000010000000001,
31'b0001110000010000000000000000000,
31'b0110100000000000000000010000100,
31'b0001110000010100000000000000000,
31'b1100000000000000000000010100001,
31'b1001000000000000010000100001000,
31'b0110000000000100000100000010000,
31'b0110000000000010000100000010000,
31'b0110000000000000000100000010000,
31'b0001110000100000000000000000000,
31'b0001000010000000001000000000010,
31'b0001110000100100000000000000000,
31'b0010000010000001000101000000000,
31'b0011000001000000000000100000010,
31'b0001010101000000000000010000000,
31'b1000001000000000000010000100001,
31'b1000000100000000000000011000001,
31'b0001110000110000000000000000000,
31'b0001010000000000100010001000000,
31'b0001000000000000100000000001010,
31'b1000000001000000100010000000001,
31'b0110000101000000000000000000100,
31'b0000000110000000000100001000000,
31'b0100000000000000100000001000001,
31'b0110000000100000000100000010000,
31'b0010000000000000000000001100100,
31'b0100100000000000000001001001000,
31'b1000100000000000000000001000001,
31'b1000100000000010000000001000001,
31'b0011000000100000000000100000010,
31'b0001100000000000000001000000011,
31'b1000100000001000000000001000001,
31'b0000110000000000000000000011000,
31'b0111000000000000000100000001000,
31'b1000000000000100010000100010000,
31'b1000100000010000000000001000001,
31'b1000000000000000010000100010000,
31'b0110000100100000000000000000100,
31'b0000001100000100000000000000001,
31'b0000001100000010000000000000001,
31'b0000001100000000000000000000001,
31'b0011000000001000000000100000010,
31'b0001010100001000000000010000000,
31'b1000100000100000000000001000001,
31'b1010000000000000000001101000000,
31'b0011000000000000000000100000010,
31'b0001010100000000000000010000000,
31'b0011000000000100000000100000010,
31'b0001010100000100000000010000000,
31'b0110000100001000000000000000100,
31'b0000000100000000011010000000000,
31'b1001100000000000000100100000000,
31'b1000000000000000100010000000001,
31'b0110000100000000000000000000100,
31'b0000000000000000100000000010010,
31'b0110000100000100000000000000100,
31'b0000001100100000000000000000001,
31'b0100000000000010000100000100000,
31'b0100000000000000000100000100000,
31'b0100010100000000000010100000000,
31'b0100000000000100000100000100000,
31'b0100010000000001100000000000001,
31'b0100000000001000000100000100000,
31'b1000001001000000010000000001000,
31'b0100100010000000000010000000001,
31'b0100010001000000000001000000100,
31'b0100000000010000000100000100000,
31'b0010001000101000000000000000010,
31'b1100000000000000000010000010100,
31'b0100001001000000100100000000000,
31'b0100000000000000000000000000111,
31'b0010001000100000000000000000010,
31'b0110000010000000000100000010000,
31'b1000101000000000000100000000000,
31'b0001000000000000001000000000010,
31'b1000101000000100000100000000000,
31'b0010000000000001000101000000000,
31'b1000101000001000000100000000000,
31'b0001000000001000001000000000010,
31'b1000000000000000001001001000000,
31'b1001001100000001000000000000000,
31'b1010000100000001001000000000000,
31'b0001000000010000001000000000010,
31'b0010001000001000000000000000010,
31'b0010001000001010000000000000010,
31'b0010001000000100000000000000010,
31'b0000000100000000000100001000000,
31'b0010001000000000000000000000010,
31'b0010001000000010000000000000010,
31'b0100010000010000000001000000100,
31'b0100000001000000000100000100000,
31'b1000100010000000000000001000001,
31'b0100000001000100000100000100000,
31'b1000001000000100010000000001000,
31'b1010000000000000010000100100000,
31'b1000001000000000010000000001000,
31'b1000010100000000000000101000000,
31'b0100010000000000000001000000100,
31'b0100010000000010000001000000100,
31'b0000111000000000000000100000000,
31'b1000010000000000000000000001101,
31'b0100001000000000100100000000000,
31'b0100001000000010100100000000000,
31'b0000000000000000000000001010100,
31'b0000001110000000000000000000001,
31'b1000101001000000000100000000000,
31'b0001000001000000001000000000010,
31'b0100000100000000000000000110100,
31'b0100000000000000001011000000000,
31'b0011000010000000000000100000010,
31'b0001010110000000000000010000000,
31'b0010000000000000010001000000100,
31'b0100100000000000010000000101000,
31'b1100000100000000000110000000000,
31'b0001000001010000001000000000010,
31'b0010010000000001000000000100100,
31'b1100010000000000000000100100000,
31'b0110000110000000000000000000100,
31'b0000000101000000000100001000000,
31'b0010001001000000000000000000010,
31'b0010001001000010000000000000010,
31'b0001110100000000000000000000000,
31'b0100100000000001100000100000000,
31'b0000000000000000100000000100001,
31'b0000010000001001000100000000000,
31'b0001110100001000000000000000000,
31'b0001000010000000000000100000001,
31'b0000010000000011000100000000000,
31'b0000010000000001000100000000000,
31'b0001110100010000000000000000000,
31'b0000001001001100000000000000001,
31'b0000011000000000000001000000010,
31'b0000001001001000000000000000001,
31'b0110000001100000000000000000100,
31'b0000001001000100000000000000001,
31'b0000001001000010000000000000001,
31'b0000001001000000000000000000001,
31'b0001110100100000000000000000000,
31'b0001010001001000000000010000000,
31'b0000010000000000000000010011000,
31'b1010000000000001100000000001000,
31'b0110000001010000000000000000100,
31'b0001010001000000000000010000000,
31'b1000000000000010000000011000001,
31'b1000000000000000000000011000001,
31'b1010000010000001001000000000000,
31'b0000000010001000000100001000000,
31'b0001100000000000000001000110000,
31'b0000101010000000001001000000000,
31'b0110000001000000000000000000100,
31'b0000000010000000000100001000000,
31'b0110000001000100000000000000100,
31'b0000001001100000000000000000001,
31'b0011000000000000001000000000001,
31'b0011000000000010001000000000001,
31'b0000010000000000010000000000100,
31'b0000010000000010010000000000100,
31'b0110000000110000000000000000100,
31'b0001010000100000000000010000000,
31'b0000010000001000010000000000100,
31'b0000001000010000000000000000001,
31'b0110000000101000000000000000100,
31'b0000001000001100000000000000001,
31'b0000010000010000010000000000100,
31'b0000001000001000000000000000001,
31'b0110000000100000000000000000100,
31'b0000001000000100000000000000001,
31'b0000001000000010000000000000001,
31'b0000001000000000000000000000001,
31'b0110000000011000000000000000100,
31'b0001010000001000000000010000000,
31'b0100000000000000000010010000001,
31'b0101001000000000001000000000100,
31'b0110000000010000000000000000100,
31'b0001010000000000000000010000000,
31'b0110000000010100000000000000100,
31'b0001010000000100000000010000000,
31'b0110000000001000000000000000100,
31'b0000000000000000011010000000000,
31'b0110000000001100000000000000100,
31'b0000001000101000000000000000001,
31'b0110000000000000000000000000100,
31'b1000000000000001000000100000000,
31'b0110000000000100000000000000100,
31'b0000001000100000000000000000001,
31'b0100010000000100000010100000000,
31'b0100000100000000000100000100000,
31'b0100010000000000000010100000000,
31'b0100010000000010000010100000000,
31'b0001000000000010000000100000001,
31'b0001000000000000000000100000001,
31'b0101100000000001000000000100000,
31'b0001000000000100000000100000001,
31'b1010000000100001001000000000000,
31'b0000000000101000000100001000000,
31'b1100000000000000001001000100000,
31'b0000101000100000001001000000000,
31'b0010000000000000100000000010001,
31'b0000000000100000000100001000000,
31'b0010001100100000000000000000010,
31'b0000001011000000000000000000001,
31'b1010000000010001001000000000000,
31'b0001000100000000001000000000010,
31'b0100010000100000000010100000000,
31'b1010100000000000000000001000010,
31'b0011100000000000000001000000000,
31'b0000000000010000000100001000000,
31'b1001001000000011000000000000000,
31'b1001001000000001000000000000000,
31'b1010000000000001001000000000000,
31'b0000000000001000000100001000000,
31'b1010000000000101001000000000000,
31'b0000101000000000001001000000000,
31'b0000000000000010000100001000000,
31'b0000000000000000000100001000000,
31'b0010001100000000000000000000010,
31'b0000000000000100000100001000000,
31'b0011000010000000001000000000001,
31'b1100000000000000000001100010000,
31'b0000010010000000010000000000100,
31'b1000101000000000000000000010100,
31'b1000001000000010000100010000000,
31'b1000001000000000000100010000000,
31'b1000010000000010000000101000000,
31'b1000010000000000000000101000000,
31'b1100000000100000000110000000000,
31'b0000101000000000000110000100000,
31'b0000111100000000000000100000000,
31'b0000100000000000010000001001000,
31'b0110000010100000000000000000100,
31'b0000001010000100000000000000001,
31'b0000001010000010000000000000001,
31'b0000001010000000000000000000001,
31'b1100000000010000000110000000000,
31'b0001010010001000000000010000000,
31'b0100000000000000000000000110100,
31'b0100000100000000001011000000000,
31'b0110000010010000000000000000100,
31'b0001010010000000000000010000000,
31'b0110100000000000000010000000010,
31'b1001001001000001000000000000000,
31'b1100000000000000000110000000000,
31'b0000000010000000011010000000000,
31'b1100000000000100000110000000000,
31'b0000101001000000001001000000000,
31'b0110000010000000000000000000100,
31'b0000000001000000000100001000000,
31'b0110000010000100000000000000100,
31'b0000001010100000000000000000001,
31'b0001111000000000000000000000000,
31'b1001000010000000010000000010000,
31'b0001111000000100000000000000000,
31'b0010000000010000000001110000000,
31'b0010100000100000000010000000100,
31'b0010000000010000100000001000100,
31'b1000000011000000010000000001000,
31'b0010000000000001000010000001000,
31'b0001111000010000000000000000000,
31'b0010000000001000100000001000100,
31'b0000100000100000000000010000001,
31'b0010000000000000000001110000000,
31'b0100000100000000000000001010010,
31'b0010000000000000100000001000100,
31'b0010000010100000000000000000010,
31'b0000000101000000000000000000001,
31'b0000000000000000000000000110010,
31'b0100100000000000011000000000000,
31'b0000100000010000000000010000001,
31'b0100100000000100011000000000000,
31'b0010100000000000000010000000100,
31'b0100100000001000011000000000000,
31'b1000000000000000000010000100001,
31'b1001000110000001000000000000000,
31'b0000100000000100000000010000001,
31'b0100100000010000011000000000000,
31'b0000100000000000000000010000001,
31'b0000100000000010000000010000001,
31'b0010000010000100000000000000010,
31'b0010000010000110000000000000010,
31'b0010000010000000000000000000010,
31'b0010000010000010000000000000010,
31'b0011000000000001000010000010000,
31'b0010000100000000000010010000100,
31'b1000101000000000000000001000001,
31'b0000000100011000000000000000001,
31'b1000000010000100010000000001000,
31'b0000000100010100000000000000001,
31'b1000000010000000010000000001000,
31'b0000000100010000000000000000001,
31'b0101010100000000000010000000000,
31'b0000000100001100000000000000001,
31'b0000110010000000000000100000000,
31'b0000000100001000000000000000001,
31'b0100000010000000100100000000000,
31'b0000000100000100000000000000001,
31'b0000000100000010000000000000001,
31'b0000000100000000000000000000001,
31'b0000100000000001000000101000000,
31'b0100100001000000011000000000000,
31'b0100000000000010000000001100001,
31'b0100000000000000000000001100001,
31'b0011001000000000000000100000010,
31'b0001011100000000000000010000000,
31'b1000000010100000010000000001000,
31'b0001000000000000000000000101010,
31'b0000100001000100000000010000001,
31'b0000000000000100001000100000010,
31'b0000100001000000000000010000001,
31'b0000000000000000001000100000010,
31'b0110001100000000000000000000100,
31'b0000001000000000100000000010010,
31'b0010000011000000000000000000010,
31'b0000000100100000000000000000001,
31'b1000100000100000000100000000000,
31'b1001000000000000010000000010000,
31'b1000100000100100000100000000000,
31'b1001000000000100010000000010000,
31'b1000100000101000000100000000000,
31'b1001000000001000010000000010000,
31'b1000000001000000010000000001000,
31'b1001000100100001000000000000000,
31'b1010000000000000110000100000000,
31'b1001000000010000010000000010000,
31'b0010000000101000000000000000010,
31'b0010000010000000000001110000000,
31'b0100000001000000100100000000000,
31'b0100001000000000000000000000111,
31'b0010000000100000000000000000010,
31'b0010000000100010000000000000010,
31'b1000100000000000000100000000000,
31'b1000100000000010000100000000000,
31'b1000100000000100000100000000000,
31'b1001000100001001000000000000000,
31'b1000100000001000000100000000000,
31'b1001000100000101000000000000000,
31'b0010000000010000000000000000010,
31'b1001000100000001000000000000000,
31'b1000100000010000000100000000000,
31'b1011000000000000000001001000000,
31'b0010000000001000000000000000010,
31'b0010000000001010000000000000010,
31'b0010000000000100000000000000010,
31'b0010000000000110000000000000010,
31'b0010000000000000000000000000010,
31'b0010000000000010000000000000010,
31'b1000100001100000000100000000000,
31'b1001000001000000010000000010000,
31'b1000000000001000010000000001000,
31'b1000100100000000000000000010100,
31'b1000000000000100010000000001000,
31'b1000000100000000000100010000000,
31'b1000000000000000010000000001000,
31'b1000000000000010010000000001000,
31'b0100000000001000100100000000000,
31'b0100010000000001000000000100001,
31'b0000110000000000000000100000000,
31'b0000110000000010000000100000000,
31'b0100000000000000100100000000000,
31'b0100000000000010100100000000000,
31'b0000000000000000001001010000000,
31'b0000000110000000000000000000001,
31'b1000100001000000000100000000000,
31'b1001000000000000000000010001100,
31'b1000100001000100000100000000000,
31'b0100001000000000001011000000000,
31'b1000100001001000000100000000000,
31'b1000100000000001010000000000100,
31'b1000000000100000010000000001000,
31'b1001000101000001000000000000000,
31'b1110010000000000000000000001000,
31'b0011000000000000000000000011010,
31'b0010000001001000000000000000010,
31'b0010010000000000000001000000001,
31'b0100000000100000100100000000000,
31'b0110000000000000000000001010001,
31'b0010000001000000000000000000010,
31'b0010000001000010000000000000010,
31'b0001111100000000000000000000000,
31'b0010000001000000000010010000100,
31'b0000010000010000000001000000010,
31'b0000000001011000000000000000001,
31'b0100000001000000011000010000000,
31'b0000000001010100000000000000001,
31'b0000000001010010000000000000001,
31'b0000000001010000000000000000001,
31'b0001000000000000000000000011001,
31'b0000000001001100000000000000001,
31'b0000010000000000000001000000010,
31'b0000000001001000000000000000001,
31'b0100000000000000000000001010010,
31'b0000000001000100000000000000001,
31'b0000000001000010000000000000001,
31'b0000000001000000000000000000001,
31'b0000100000000000100001000001000,
31'b0110000000000000100000000100100,
31'b0000100100010000000000010000001,
31'b1100100000000000100000000000001,
31'b0110000000000000010001000000010,
31'b1001000010000101000000000000000,
31'b1001000010000011000000000000000,
31'b1001000010000001000000000000000,
31'b0001010000000000100000010100000,
31'b0000100010000100001001000000000,
31'b0000100100000000000000010000001,
31'b0000100010000000001001000000000,
31'b0110001001000000000000000000100,
31'b0000001010000000000100001000000,
31'b0010000110000000000000000000010,
31'b0000000001100000000000000000001,
31'b0101010000010000000010000000000,
31'b0010000000000000000010010000100,
31'b0000011000000000010000000000100,
31'b0000000000011000000000000000001,
31'b0100000000000000011000010000000,
31'b0000000000010100000000000000001,
31'b0000000000010010000000000000001,
31'b0000000000010000000000000000001,
31'b0101010000000000000010000000000,
31'b0000000000001100000000000000001,
31'b0000000000001010000000000000001,
31'b0000000000001000000000000000001,
31'b0000000000000110000000000000001,
31'b0000000000000100000000000000001,
31'b0000000000000010000000000000001,
31'b0000000000000000000000000000001,
31'b1000000010000001000000000011000,
31'b0110010000000000010000000000001,
31'b0101000000000010001000000000100,
31'b0101000000000000001000000000100,
31'b0110001000010000000000000000100,
31'b0001011000000000000000010000000,
31'b0011000000000000010010000000000,
31'b0000000000110000000000000000001,
31'b0110001000001000000000000000100,
31'b0000001000000000011010000000000,
31'b0010010000000000001000010000000,
31'b0000000000101000000000000000001,
31'b0110001000000000000000000000100,
31'b0000000000100100000000000000001,
31'b0000000000100010000000000000001,
31'b0000000000100000000000000000001,
31'b1000100100100000000100000000000,
31'b1001000100000000010000000010000,
31'b0110000000000000000000001100010,
31'b1001000000101001000000000000000,
31'b1001100000000000000000000001100,
31'b1000000001000000000100010000000,
31'b1001000000100011000000000000000,
31'b1001000000100001000000000000000,
31'b0010000000000100001000100000001,
31'b0000100001000000000110000100000,
31'b0010000000000000001000100000001,
31'b0000100000100000001001000000000,
31'b0100000101000000100100000000000,
31'b0000001000100000000100001000000,
31'b0010000100100000000000000000010,
31'b0000000011000000000000000000001,
31'b1000100100000000000100000000000,
31'b1001000000001101000000000000000,
31'b1001000000001011000000000000000,
31'b1001000000001001000000000000000,
31'b1001000000000111000000000000000,
31'b1001000000000101000000000000000,
31'b1001000000000011000000000000000,
31'b1001000000000001000000000000000,
31'b1010001000000001001000000000000,
31'b0000100000000100001001000000000,
31'b0010000100001000000000000000010,
31'b0000100000000000001001000000000,
31'b0010000100000100000000000000010,
31'b0000001000000000000100001000000,
31'b0010000100000000000000000000010,
31'b0000010000000000000000110000000,
31'b1000000000100001000000000011000,
31'b1000000000001000000100010000000,
31'b1000100000000010000000000010100,
31'b1000100000000000000000000010100,
31'b1000000000000010000100010000000,
31'b1000000000000000000100010000000,
31'b1000000100000000010000000001000,
31'b0000000010010000000000000000001,
31'b0101010010000000000010000000000,
31'b0000100000000000000110000100000,
31'b0000110100000000000000100000000,
31'b0000000010001000000000000000001,
31'b0100000100000000100100000000000,
31'b0000000010000100000000000000001,
31'b0000000010000010000000000000001,
31'b0000000010000000000000000000001,
31'b1000000000000001000000000011000,
31'b1000000000101000000100010000000,
31'b1001000000000000010100000000100,
31'b1001000001001001000000000000000,
31'b1000000000100010000100010000000,
31'b1000000000100000000100010000000,
31'b1001000001000011000000000000000,
31'b1001000001000001000000000000000,
31'b1100001000000000000110000000000,
31'b0000100001000100001001000000000,
31'b0010010010000000001000010000000,
31'b0000100001000000001001000000000,
31'b0110001010000000000000000000100,
31'b0000001001000000000100001000000,
31'b0010000101000000000000000000010,
31'b0000000010100000000000000000001,
31'b0010000000000000000000000000000,
31'b0010000000000010000000000000000,
31'b0010000000000100000000000000000,
31'b0010000000000110000000000000000,
31'b0010000000001000000000000000000,
31'b0010000000001010000000000000000,
31'b0010000000001100000000000000000,
31'b0010000000001110000000000000000,
31'b0010000000010000000000000000000,
31'b0010000000010010000000000000000,
31'b0010000000010100000000000000000,
31'b0010000000010110000000000000000,
31'b0010000000011000000000000000000,
31'b0010000000011010000000000000000,
31'b0000000010000000000000000110000,
31'b0001001000000000001000000000000,
31'b0010000000100000000000000000000,
31'b0010000000100010000000000000000,
31'b0010000000100100000000000000000,
31'b0100001000000000000000000000101,
31'b0010000000101000000000000000000,
31'b0010000000101010000000000000000,
31'b0100010000010000010000000000000,
31'b0100010000010010010000000000000,
31'b0010000000110000000000000000000,
31'b0010000000110010000000000000000,
31'b0100010000001000010000000000000,
31'b0100010000001010010000000000000,
31'b0100010000000100010000000000000,
31'b0110001000000000000010010000000,
31'b0100010000000000010000000000000,
31'b0100010000000010010000000000000,
31'b0010000001000000000000000000000,
31'b0010000001000010000000000000000,
31'b0010000001000100000000000000000,
31'b0010000001000110000000000000000,
31'b0010000001001000000000000000000,
31'b0000000010000000001000100000000,
31'b0010000001001100000000000000000,
31'b0011000000000000000000000011000,
31'b0010000001010000000000000000000,
31'b0010000001010010000000000000000,
31'b0010000001010100000000000000000,
31'b0010000001010110000000000000000,
31'b0010000001011000000000000000000,
31'b0010001000000000100000000100000,
31'b0000000000000000100000100001000,
31'b0001001001000000001000000000000,
31'b0010000001100000000000000000000,
31'b0010000001100010000000000000000,
31'b0100000000000000100100000000010,
31'b0100001001000000000000000000101,
31'b0010000001101000000000000000000,
31'b0010100100000000000000010000000,
31'b0100010001010000010000000000000,
31'b1001000000000000001000011000000,
31'b1000000000000000010000000001010,
31'b1010000100000000000010000100000,
31'b1010010000000000000100100000000,
31'b1000010000000000010010001000000,
31'b1110100000000000100000000000000,
31'b0010100100010000000000010000000,
31'b0100010001000000010000000000000,
31'b0100010001000010010000000000000,
31'b0010000010000000000000000000000,
31'b0010000010000010000000000000000,
31'b0010000010000100000000000000000,
31'b0010000010000110000000000000000,
31'b0010000010001000000000000000000,
31'b0000000001000000001000100000000,
31'b0000000000010000000000000110000,
31'b0000000001000100001000100000000,
31'b0010000010010000000000000000000,
31'b0010000010010010000000000000000,
31'b0000000000001000000000000110000,
31'b0010000000000000101000000001000,
31'b0000000000000100000000000110000,
31'b0000000001010000001000100000000,
31'b0000000000000000000000000110000,
31'b0000000000000010000000000110000,
31'b0010000010100000000000000000000,
31'b0010000010100010000000000000000,
31'b0100000100000000000000001010000,
31'b0100001010000000000000000000101,
31'b0000010100000000000001000000000,
31'b0000010100000010000001000000000,
31'b0000010100000100000001000000000,
31'b1000010000010000001100000000000,
31'b0010000010110000000000000000000,
31'b0010000010110010000000000000000,
31'b0010010000000001000000001000000,
31'b1000010000001000001100000000000,
31'b0000010100010000000001000000000,
31'b1000010000000100001100000000000,
31'b0000000000100000000000000110000,
31'b1000010000000000001100000000000,
31'b0010000011000000000000000000000,
31'b0000000000001000001000100000000,
31'b0010000011000100000000000000000,
31'b0000001000000000100000000010000,
31'b0000000000000010001000100000000,
31'b0000000000000000001000100000000,
31'b0000000001010000000000000110000,
31'b0000000000000100001000100000000,
31'b0010000011010000000000000000000,
31'b0001000000000000000000000101000,
31'b0011001000000000000000100000000,
31'b0001000000000100000000000101000,
31'b0000000001000100000000000110000,
31'b0000000000010000001000100000000,
31'b0000000001000000000000000110000,
31'b0000000001000010000000000110000,
31'b0010000011100000000000000000000,
31'b0000000100000000000000000000011,
31'b0100000101000000000000001010000,
31'b0000001000100000100000000010000,
31'b0000010101000000000001000000000,
31'b0000000000100000001000100000000,
31'b1000000100000010000010000010000,
31'b1000000100000000000010000010000,
31'b1011000000000001000000000000001,
31'b0001000000100000000000000101000,
31'b0011001000100000000000100000000,
31'b0001101000000000000001000000001,
31'b0000010101010000000001000000000,
31'b0000000100000000000100000100100,
31'b0000010000000000000010100000100,
31'b1000010001000000001100000000000,
31'b0010000100000000000000000000000,
31'b0010000100000010000000000000000,
31'b0010000100000100000000000000000,
31'b0010000100000110000000000000000,
31'b0010000100001000000000000000000,
31'b0010000100001010000000000000000,
31'b0010000100001100000000000000000,
31'b0011100000000001000100000000000,
31'b0010000100010000000000000000000,
31'b1001000000000001000000000000010,
31'b0010000100010100000000000000000,
31'b1010000000000000001101000000000,
31'b0010000100011000000000000000000,
31'b1010101000000000000000001000000,
31'b0000000000000001000001001000000,
31'b0001001100000000001000000000000,
31'b0010000100100000000000000000000,
31'b0010000100100010000000000000000,
31'b0100000010000000000000001010000,
31'b0100001100000000000000000000101,
31'b0000010010000000000001000000000,
31'b0010100001000000000000010000000,
31'b0010000000000001010000000010000,
31'b1000010000000000110000010000000,
31'b0010000100110000000000000000000,
31'b1010000001000000000010000100000,
31'b0100010100001000010000000000000,
31'b1001000000000000101010000000000,
31'b0110000000000000000000001100000,
31'b0110000000000010000000001100000,
31'b0100010100000000010000000000000,
31'b0100010100000010010000000000000,
31'b0010000101000000000000000000000,
31'b0010000101000010000000000000000,
31'b0010000101000100000000000000000,
31'b0010000101000110000000000000000,
31'b0010000101001000000000000000000,
31'b0010100000100000000000010000000,
31'b0010000101001100000000000000000,
31'b1100000000000000000000110001000,
31'b0010000101010000000000000000000,
31'b1010000000100000000010000100000,
31'b0010000101010100000000000000000,
31'b1100000000000001000011000000000,
31'b0010000101011000000000000000000,
31'b0010100000110000000000010000000,
31'b0000000100000000100000100001000,
31'b0101010000000001000000000001000,
31'b0010000101100000000000000000000,
31'b0000000010000000000000000000011,
31'b0100000100000000100100000000010,
31'b0010000000000000000100000010100,
31'b0010100000000010000000010000000,
31'b0010100000000000000000010000000,
31'b1000001000000001000001010000000,
31'b1000000010000000000010000010000,
31'b1010000000000010000010000100000,
31'b1010000000000000000010000100000,
31'b1000001000000000000010100001000,
31'b1000000000000000000100010000010,
31'b0110000001000000000000001100000,
31'b0010100000010000000000010000000,
31'b0101000000000000101000001000000,
31'b1000000010010000000010000010000,
31'b0010000110000000000000000000000,
31'b0010000110000010000000000000000,
31'b0100000000100000000000001010000,
31'b0110000000000000100100000000001,
31'b0000010000100000000001000000000,
31'b0000010000100010000001000000000,
31'b0000010000100100000001000000000,
31'b1000010000000000000000100100100,
31'b0010000110010000000000000000000,
31'b1010000000000000010000000001001,
31'b0110000000000000010001000000000,
31'b0110000000000010010001000000000,
31'b0000010000110000000001000000000,
31'b0000010000110010000001000000000,
31'b0000000100000000000000000110000,
31'b0000000100000010000000000110000,
31'b0000010000001000000001000000000,
31'b0000000001000000000000000000011,
31'b0100000000000000000000001010000,
31'b0100000000000010000000001010000,
31'b0000010000000000000001000000000,
31'b0000010000000010000001000000000,
31'b0000010000000100000001000000000,
31'b1000000001000000000010000010000,
31'b0000000000000001010000000100000,
31'b0000000001010000000000000000011,
31'b0100000000010000000000001010000,
31'b0100100000000000010000100000001,
31'b0000010000010000000001000000000,
31'b0000010000010010000001000000000,
31'b0000010000010100000001000000000,
31'b1000010100000000001100000000000,
31'b0010000111000000000000000000000,
31'b0000000000100000000000000000011,
31'b0110001000000000000000000000110,
31'b0000001100000000100000000010000,
31'b0000010001100000000001000000000,
31'b0000000100000000001000100000000,
31'b1000000000100010000010000010000,
31'b1000000000100000000010000010000,
31'b0011000000000000010010000000010,
31'b0001000100000000000000000101000,
31'b1100001000000000000000010010000,
31'b0001011000000000000000010000010,
31'b1000010000000000001000000010100,
31'b0000000100010000001000100000000,
31'b1000000000000000000101100000000,
31'b1000000000110000000010000010000,
31'b0000000000000010000000000000011,
31'b0000000000000000000000000000011,
31'b0100000001000000000000001010000,
31'b0000000000000100000000000000011,
31'b0000010001000000000001000000000,
31'b0000000000001000000000000000011,
31'b1000000000000010000010000010000,
31'b1000000000000000000010000010000,
31'b0000000001000001010000000100000,
31'b0000000000010000000000000000011,
31'b0100000001010000000000001010000,
31'b0000100000000000000000010110000,
31'b0000010001010000000001000000000,
31'b0000000000000000000100000100100,
31'b1000000000100000000101100000000,
31'b1000000000010000000010000010000,
31'b0010001000000000000000000000000,
31'b0010001000000010000000000000000,
31'b0010001000000100000000000000000,
31'b0000000000000000000000100101000,
31'b0010001000001000000000000000000,
31'b0010001000001010000000000000000,
31'b0010001000001100000000000000000,
31'b0001000000010000001000000000000,
31'b0010001000010000000000000000000,
31'b0010001000010010000000000000000,
31'b0010001000010100000000000000000,
31'b0001000000001000001000000000000,
31'b0010001000011000000000000000000,
31'b0001000000000100001000000000000,
31'b0001000000000010001000000000000,
31'b0001000000000000001000000000000,
31'b0010001000100000000000000000000,
31'b0100000000000100000000000000101,
31'b0100000000000010000000000000101,
31'b0100000000000000000000000000101,
31'b0010001000101000000000000000000,
31'b0110000000010000000010010000000,
31'b0100011000010000010000000000000,
31'b0100000000001000000000000000101,
31'b0010001000110000000000000000000,
31'b0110000000001000000010010000000,
31'b0100011000001000010000000000000,
31'b0100000000010000000000000000101,
31'b0110000000000010000010010000000,
31'b0110000000000000000010010000000,
31'b0100011000000000010000000000000,
31'b0001000000100000001000000000000,
31'b0010001001000000000000000000000,
31'b0010001001000010000000000000000,
31'b0010001001000100000000000000000,
31'b0000000010000000100000000010000,
31'b0010001001001000000000000000000,
31'b0010000000010000100000000100000,
31'b0010001001001100000000000000000,
31'b0001000001010000001000000000000,
31'b0000000000000000001000000011000,
31'b0010000000001000100000000100000,
31'b0011000010000000000000100000000,
31'b0001000001001000001000000000000,
31'b0010000000000010100000000100000,
31'b0010000000000000100000000100000,
31'b0001000001000010001000000000000,
31'b0001000001000000001000000000000,
31'b0010001001100000000000000000000,
31'b0110000100000000100000001000000,
31'b0100001000000000100100000000010,
31'b0100000001000000000000000000101,
31'b0010100000000000000010001100000,
31'b0010101100000000000000010000000,
31'b1000000100000001000001010000000,
31'b1001000000000000000001000010100,
31'b1010000000000000000000011000000,
31'b1010000000000010000000011000000,
31'b1010000000000100000000011000000,
31'b0100000001010000000000000000101,
31'b1010000000001000000000011000000,
31'b0010000000100000100000000100000,
31'b0100011001000000010000000000000,
31'b0100000000000001100001000000000,
31'b0010001010000000000000000000000,
31'b0010001010000010000000000000000,
31'b0010001010000100000000000000000,
31'b0000000001000000100000000010000,
31'b0001000000000000100000000001000,
31'b0001000000000010100000000001000,
31'b0001000000000100100000000001000,
31'b0001000010010000001000000000000,
31'b0010001010010000000000000000000,
31'b0010001010010010000000000000000,
31'b0011000001000000000000100000000,
31'b0001000010001000001000000000000,
31'b0001000000010000100000000001000,
31'b0010000000000000000000100011000,
31'b0000001000000000000000000110000,
31'b0001000010000000001000000000000,
31'b0010001010100000000000000000000,
31'b0110000000000000000100000010010,
31'b0100001100000000000000001010000,
31'b0100000010000000000000000000101,
31'b0001000000100000100000000001000,
31'b0001010000000001001000001000000,
31'b0001110000010000000000000000010,
31'b1100100000010000000000000010000,
31'b0010001010110000000000000000000,
31'b1100000000000000000100010000100,
31'b0011000001100000000000100000000,
31'b1100100000001000000000000010000,
31'b0001110000000100000000000000010,
31'b1100100000000100000000000010000,
31'b0001110000000000000000000000010,
31'b1100100000000000000000000010000,
31'b0010001011000000000000000000000,
31'b0000000000000100100000000010000,
31'b0000000000000010100000000010000,
31'b0000000000000000100000000010000,
31'b0001000001000000100000000001000,
31'b0000001000000000001000100000000,
31'b0010000000000000001000000101000,
31'b0000000000001000100000000010000,
31'b0011000000000100000000100000000,
31'b0001001000000000000000000101000,
31'b0011000000000000000000100000000,
31'b0000000000010000100000000010000,
31'b0011000000001100000000100000000,
31'b0010000010000000100000000100000,
31'b0011000000001000000000100000000,
31'b0001000011000000001000000000000,
31'b0010001011100000000000000000000,
31'b0000001100000000000000000000011,
31'b0010000000000000000100001000001,
31'b0000000000100000100000000010000,
31'b0101010000000000010000100000000,
31'b0000001000100000001000100000000,
31'b1000000000000011001000000000001,
31'b1000000000000001001000000000001,
31'b1101100000000000000000000001000,
31'b0001100000000100000001000000001,
31'b0011000000100000000000100000000,
31'b0001100000000000000001000000001,
31'b1100000000000001010000010000000,
31'b0010000010100000100000000100000,
31'b0011000000101000000000100000000,
31'b1100100001000000000000000010000,
31'b0010001100000000000000000000000,
31'b0010001100000010000000000000000,
31'b0010001100000100000000000000000,
31'b0000000000000000000100001000010,
31'b1001000000000000000101000000000,
31'b1010100000010000000000001000000,
31'b1010000000000001001000000000010,
31'b0001000100010000001000000000000,
31'b0010001100010000000000000000000,
31'b1010100000001000000000001000000,
31'b0011100000000000000001000000010,
31'b0001000100001000001000000000000,
31'b1010100000000010000000001000000,
31'b1010100000000000000000001000000,
31'b0001000100000010001000000000000,
31'b0001000100000000001000000000000,
31'b0010001100100000000000000000000,
31'b0110000001000000100000001000000,
31'b0100001010000000000000001010000,
31'b0100000100000000000000000000101,
31'b1010000000000000100010000000000,
31'b1010000000000010100010000000000,
31'b1010000000000100100010000000000,
31'b0100000100001000000000000000101,
31'b0010100000000000100000010100000,
31'b0001000000000100000000100000011,
31'b1000000001000000000010100001000,
31'b0001000000000000000000100000011,
31'b1010000000010000100010000000000,
31'b1010100000100000000000001000000,
31'b0100011100000000010000000000000,
31'b0100000000000000000000101001000,
31'b0100000000000000000100000010001,
31'b0110000000100000100000001000000,
31'b0110000010000000000000000000110,
31'b0000000110000000100000000010000,
31'b1110000000000000000000010100000,
31'b0010101000100000000000010000000,
31'b1100000000000000000110000000010,
31'b0001010000000000000110000010000,
31'b0110100000000000000010000000000,
31'b0110100000000010000010000000000,
31'b1100000010000000000000010010000,
31'b0001010010000000000000010000010,
31'b0110100000001000000010000000000,
31'b0010000100000000100000000100000,
31'b0001010000100000000001100000000,
31'b0001000101000000001000000000000,
31'b0110000000000010100000001000000,
31'b0110000000000000100000001000000,
31'b1000000000010000000010100001000,
31'b0110000000000100100000001000000,
31'b1010000001000000100010000000000,
31'b0010101000000000000000010000000,
31'b1000000000000001000001010000000,
31'b1000001010000000000010000010000,
31'b1010000100000000000000011000000,
31'b1010001000000000000010000100000,
31'b1000000000000000000010100001000,
31'b1000001000000000000100010000010,
31'b0001010000000100000001100000000,
31'b0010101000010000000000010000000,
31'b0001010000000000000001100000000,
31'b0100000100000001100001000000000,
31'b0010001110000000000000000000000,
31'b0010001110000010000000000000000,
31'b0110000001000000000000000000110,
31'b0000000101000000100000000010000,
31'b0001000100000000100000000001000,
31'b0101000000000000011001000000000,
31'b0001000100000100100000000001000,
31'b0001000110010000001000000000000,
31'b0010100000000000010000100000100,
31'b1100100000000001010000000000000,
31'b1100000001000000000000010010000,
31'b0001010001000000000000010000010,
31'b0001000100010000100000000001000,
31'b1101000000000000000000010001000,
31'b0001000000000000000001010000001,
31'b0001000110000000001000000000000,
31'b0000000000000000100100000000100,
31'b0000001001000000000000000000011,
31'b0100001000000000000000001010000,
31'b0100001000000010000000001010000,
31'b0000011000000000000001000000000,
31'b0000011000000010000001000000000,
31'b0000100000000000100000010010000,
31'b1010110000000001000000000000000,
31'b0000001000000001010000000100000,
31'b0000010000000001000100000000010,
31'b1100000000000000010000000001100,
31'b0011010000000000001001000000000,
31'b0000011000010000000001000000000,
31'b0000011000010010000001000000000,
31'b0001110100000000000000000000010,
31'b1100100100000000000000000010000,
31'b0110000000000100000000000000110,
31'b0000001000100000000000000000011,
31'b0110000000000000000000000000110,
31'b0000000100000000100000000010000,
31'b0001000101000000100000000001000,
31'b0000001100000000001000100000000,
31'b0110000000001000000000000000110,
31'b0000000100001000100000000010000,
31'b1100000000000100000000010010000,
31'b0001010000000100000000010000010,
31'b1100000000000000000000010010000,
31'b0001010000000000000000010000010,
31'b1100100000000000000100000000100,
31'b0010100000000001000100100000000,
31'b1100000000001000000000010010000,
31'b0001010000001000000000010000010,
31'b0000001000000010000000000000011,
31'b0000001000000000000000000000011,
31'b0110000000100000000000000000110,
31'b0000001000000100000000000000011,
31'b0000011001000000000001000000000,
31'b0000000000000001110000000000000,
31'b1000001000000010000010000010000,
31'b1000001000000000000010000010000,
31'b0000010000001000010000000000110,
31'b0000010000000000100001000100000,
31'b1100000000100000000000010010000,
31'b0001100100000000000001000000001,
31'b0000010000000000010000000000110,
31'b0000001000000000000100000100100,
31'b0011000000000000001000000000011,
31'b1100000000000001000100000001000,
31'b0010010000000000000000000000000,
31'b0010010000000010000000000000000,
31'b0010010000000100000000000000000,
31'b0010010000000110000000000000000,
31'b0010010000001000000000000000000,
31'b0010010000001010000000000000000,
31'b0100000000110000010000000000000,
31'b0111000000000000000010000000001,
31'b0010010000010000000000000000000,
31'b0101000000000000000000010000100,
31'b0100000000101000010000000000000,
31'b0101000000000100000000010000100,
31'b0100000000100100010000000000000,
31'b0101000000001000000000010000100,
31'b0100000000100000010000000000000,
31'b0100000000100010010000000000000,
31'b0010010000100000000000000000000,
31'b0010010000100010000000000000000,
31'b0100000000011000010000000000000,
31'b0100011000000000000000000000101,
31'b0000000110000000000001000000000,
31'b0000000000000000001000010000001,
31'b0100000000010000010000000000000,
31'b0100000000010010010000000000000,
31'b0100000000001100010000000000000,
31'b0101000000100000000000010000100,
31'b0100000000001000010000000000000,
31'b0100000000001010010000000000000,
31'b0100000000000100010000000000000,
31'b0100000000000110010000000000000,
31'b0100000000000000010000000000000,
31'b0100000000000010010000000000000,
31'b0010010001000000000000000000000,
31'b0010010001000010000000000000000,
31'b1000100000000000110000000000000,
31'b1010000000000000000011000010000,
31'b0010010001001000000000000000000,
31'b0010000000000000000001000000011,
31'b1110000000000000000000000001010,
31'b0011010000000000000000000011000,
31'b0100100000000000000100000001000,
31'b0101000001000000000000010000100,
31'b1010000000100000000100100000000,
31'b1000100000000000000101000000001,
31'b0100100000001000000100000001000,
31'b1000001000000000001000001000001,
31'b0100000001100000010000000000000,
31'b0101000100000001000000000001000,
31'b0010010001100000000000000000000,
31'b0010010001100010000000000000000,
31'b1010000000010000000100100000000,
31'b1001000000000000100100000010000,
31'b0000100000000000000000100000010,
31'b0000100000000010000000100000010,
31'b0100000001010000010000000000000,
31'b0100000001010010010000000000000,
31'b1010000000000100000100100000000,
31'b1000001000000000000100000101000,
31'b1010000000000000000100100000000,
31'b1000000000000000010010001000000,
31'b0100000001000100010000000000000,
31'b0100100000000001000000010010000,
31'b0100000001000000010000000000000,
31'b0100000001000010010000000000000,
31'b0010010010000000000000000000000,
31'b0010010010000010000000000000000,
31'b0010010010000100000000000000000,
31'b0010100000000001100010000000000,
31'b0000000100100000000001000000000,
31'b0000010001000000001000100000000,
31'b0000010000010000000000000110000,
31'b1000000100000000000000100100100,
31'b0100000000000000000001001100000,
31'b0101000010000000000000010000100,
31'b0010000000100001000000001000000,
31'b1000000000101000001100000000000,
31'b0000010000000100000000000110000,
31'b1000000001000000000011000100000,
31'b0000010000000000000000000110000,
31'b1000000000100000001100000000000,
31'b0000000100001000000001000000000,
31'b0010100000000000001000000000010,
31'b0010000000010001000000001000000,
31'b1001000100000000000000001000010,
31'b0000000100000000000001000000000,
31'b0000000100000010000001000000000,
31'b0000000100000100000001000000000,
31'b1000000000010000001100000000000,
31'b0010000000000101000000001000000,
31'b1000101000000000000001001000000,
31'b0010000000000001000000001000000,
31'b1000000000001000001100000000000,
31'b0000000100010000000001000000000,
31'b1000000000000100001100000000000,
31'b0100000010000000010000000000000,
31'b1000000000000000001100000000000,
31'b0010010011000000000000000000000,
31'b0000100000000000000001010000000,
31'b1010001000000001000000010000000,
31'b0000100000000100000001010000000,
31'b0000010000000010001000100000000,
31'b0000010000000000001000100000000,
31'b0000010001010000000000000110000,
31'b0000010000000100001000100000000,
31'b0100100010000000000100000001000,
31'b0001010000000000000000000101000,
31'b0011011000000000000000100000000,
31'b0001010000000100000000000101000,
31'b1000000100000000001000000010100,
31'b1000000000000000000011000100000,
31'b0000010001000000000000000110000,
31'b1000000001100000001100000000000,
31'b0010000000000000000000110000001,
31'b0000100000100000000001010000000,
31'b0010000001010001000000001000000,
31'b0001100000000000100000000100010,
31'b0000000101000000000001000000000,
31'b0000010000100000001000100000000,
31'b0000000101000100000001000000000,
31'b1000010100000000000010000010000,
31'b0010000001000101000000001000000,
31'b0001010000100000000000000101000,
31'b0010000001000001000000001000000,
31'b1000000010000000010010001000000,
31'b0000000101010000000001000000000,
31'b1000000001000100001100000000000,
31'b0000000000000000000010100000100,
31'b1000000001000000001100000000000,
31'b0010010100000000000000000000000,
31'b0000000000000000000000110000010,
31'b0000000000000000010000001100000,
31'b0000000000000100000000110000010,
31'b0000000010100000000001000000000,
31'b0000000010100010000001000000000,
31'b0000000010100100000001000000000,
31'b1000000010000000000000100100100,
31'b0100000000000001000000000010000,
31'b0100000000000011000000000010000,
31'b0100000000000101000000000010000,
31'b0100100001000000010000010000000,
31'b0100000000001001000000000010000,
31'b0100000000100000000100010001000,
31'b0100000100100000010000000000000,
31'b0101000001000001000000000001000,
31'b0000000010001000000001000000000,
31'b0000000010001010000001000000000,
31'b0000000010001100000001000000000,
31'b1001000010000000000000001000010,
31'b0000000010000000000001000000000,
31'b0000000010000010000001000000000,
31'b0000000010000100000001000000000,
31'b1000000000000000110000010000000,
31'b0100000000100001000000000010000,
31'b0100000000100011000000000010000,
31'b0100000100001000010000000000000,
31'b0100100000000000000000000011100,
31'b0000000010010000000001000000000,
31'b0100000000000000000100010001000,
31'b0100000100000000010000000000000,
31'b0100000100000010010000000000000,
31'b0000100000000000001000000000001,
31'b0000100000000010001000000000001,
31'b0000100000000100001000000000001,
31'b0100100000010000010000010000000,
31'b0000100000001000001000000000001,
31'b0010110000100000000000010000000,
31'b0000101000100000010010000000000,
31'b1100000000000000010010000100000,
31'b0100000001000001000000000010000,
31'b0100100000000100010000010000000,
31'b0100100000000010010000010000000,
31'b0100100000000000010000010000000,
31'b1001000000000001000001000000001,
31'b1001001000000000000000000100100,
31'b0101000000000011000000000001000,
31'b0101000000000001000000000001000,
31'b0000100000100000001000000000001,
31'b0010000000000000001001100000000,
31'b0000101000001000010010000000000,
31'b0010010000000000000100000010100,
31'b0000000011000000000001000000000,
31'b0010110000000000000000010000000,
31'b0000101000000000010010000000000,
31'b1000010010000000000010000010000,
31'b0101100000001000000000000000100,
31'b1010010000000000000010000100000,
31'b1010000100000000000100100000000,
31'b1000010000000000000100010000010,
31'b0101100000000000000000000000100,
31'b0101100000000010000000000000100,
31'b0100000101000000010000000000000,
31'b0101000000100001000000000001000,
31'b0000000000101000000001000000000,
31'b0000000010000000000000110000010,
31'b0000000010000000010000001100000,
31'b1001000000100000000000001000010,
31'b0000000000100000000001000000000,
31'b0000000000100010000001000000000,
31'b0000000000100100000001000000000,
31'b1000000000000000000000100100100,
31'b0100000010000001000000000010000,
31'b0100001000000000000011010000000,
31'b0110010000000000010001000000000,
31'b1001000000000000001000000001100,
31'b0000000000110000000001000000000,
31'b0000000000110010000001000000000,
31'b0000010100000000000000000110000,
31'b1000000100100000001100000000000,
31'b0000000000001000000001000000000,
31'b0000000000001010000001000000000,
31'b0000000000001100000001000000000,
31'b1001000000000000000000001000010,
31'b0000000000000000000001000000000,
31'b0000000000000010000001000000000,
31'b0000000000000100000001000000000,
31'b0000000000000110000001000000000,
31'b0000000000011000000001000000000,
31'b0000001000000001000100000000010,
31'b0010000100000001000000001000000,
31'b1001000000010000000000001000010,
31'b0000000000010000000001000000000,
31'b0000000000010010000001000000000,
31'b0000000000010100000001000000000,
31'b1000000100000000001100000000000,
31'b0000100010000000001000000000001,
31'b0000100100000000000001010000000,
31'b0000100010000100001000000000001,
31'b0001001000010000000000010000010,
31'b0000000001100000000001000000000,
31'b0000010100000000001000100000000,
31'b0000000001100100000001000000000,
31'b1000010000100000000010000010000,
31'b1100100000000000100001000000000,
31'b0001010100000000000000000101000,
31'b1000100000000000001100010000000,
31'b0001001000000000000000010000010,
31'b1000000000000000001000000010100,
31'b1000000100000000000011000100000,
31'b1000010000000000000101100000000,
31'b0110000000000000010000000000011,
31'b0000000001001000000001000000000,
31'b0000010000000000000000000000011,
31'b0000000001001100000001000000000,
31'b0001000000000000000001000011000,
31'b0000000001000000000001000000000,
31'b0000000001000010000001000000000,
31'b0000000001000100000001000000000,
31'b1000010000000000000010000010000,
31'b0000000001011000000001000000000,
31'b0000010000010000000000000000011,
31'b0010000101000001000000001000000,
31'b0001001000100000000000010000010,
31'b0000000001010000000001000000000,
31'b0000010000000000000100000100100,
31'b0000000100000000000010100000100,
31'b1000010000010000000010000010000,
31'b0010011000000000000000000000000,
31'b0010011000000010000000000000000,
31'b0010011000000100000000000000000,
31'b0000000000000000010010010000000,
31'b0010011000001000000000000000000,
31'b0010011000001010000000000000000,
31'b0110000000000000001000010000100,
31'b0001010000010000001000000000000,
31'b0100000000000000001010000000001,
31'b0101001000000000000000010000100,
31'b0100001000101000010000000000000,
31'b0001010000001000001000000000000,
31'b0100001000100100010000000000000,
31'b0010000000000000010000000000101,
31'b0100001000100000010000000000000,
31'b0001010000000000001000000000000,
31'b0010011000100000000000000000000,
31'b0111000000000000011000000000000,
31'b0100010000000010000000000000101,
31'b0100010000000000000000000000101,
31'b0001000000000000000010000000100,
31'b0001000000000010000010000000100,
31'b0100001000010000010000000000000,
31'b0100010000001000000000000000101,
31'b0100001000001100010000000000000,
31'b1000100010000000000001001000000,
31'b0100001000001000010000000000000,
31'b0100010000010000000000000000101,
31'b0100001000000100010000000000000,
31'b0110010000000000000010010000000,
31'b0100001000000000010000000000000,
31'b0100001000000010010000000000000,
31'b0010011001000000000000000000000,
31'b0010011001000010000000000000000,
31'b1010000010000001000000010000000,
31'b0000010010000000100000000010000,
31'b0010011001001000000000000000000,
31'b1100000000000000000000100100010,
31'b1100000000000000010000011000000,
31'b0001010001010000001000000000000,
31'b0010000000000001000100000000001,
31'b1000000000100000000100000101000,
31'b0011010010000000000000100000000,
31'b0001010001001000001000000000000,
31'b1000000000000010001000001000001,
31'b1000000000000000001000001000001,
31'b0100001001100000010000000000000,
31'b0001010001000000001000000000000,
31'b0011000000000001000000101000000,
31'b1101000000000000000000001000100,
31'b0100000000001000000001000000110,
31'b0100000000000000110000000100000,
31'b0001000001000000000010000000100,
31'b1001000000000000001100100000000,
31'b0100000000000000000001000000110,
31'b0100000000001000110000000100000,
31'b1010010000000000000000011000000,
31'b1000000000000000000100000101000,
31'b1010001000000000000100100000000,
31'b1000001000000000010010001000000,
31'b0100100010000000000011000000000,
31'b1000000000100000001000001000001,
31'b0100001001000000010000000000000,
31'b0100010000000001100001000000000,
31'b1000000000000000100011000000000,
31'b1010100000000000010000000010000,
31'b1010000001000001000000010000000,
31'b0000010001000000100000000010000,
31'b0001010000000000100000000001000,
31'b0100000100000001000000100001000,
31'b0001100000110000000000000000010,
31'b0001010010010000001000000000000,
31'b1010000000000000000000101000001,
31'b1000100000100000000001001000000,
31'b0011010001000000000000100000000,
31'b0001010010001000001000000000000,
31'b0001100000100100000000000000010,
31'b0010010000000000000000100011000,
31'b0001100000100000000000000000010,
31'b0001010010000000001000000000000,
31'b1011000000000000000100000000000,
31'b1011000000000010000100000000000,
31'b1011000000000100000100000000000,
31'b0100010010000000000000000000101,
31'b0000001100000000000001000000000,
31'b0001000000000001001000001000000,
31'b0001100000010000000000000000010,
31'b1010100100000001000000000000000,
31'b1011000000010000000100000000000,
31'b1000100000000000000001001000000,
31'b0010001000000001000000001000000,
31'b1000100000000100000001001000000,
31'b0001100000000100000000000000010,
31'b1000100000001000000001001000000,
31'b0001100000000000000000000000010,
31'b1000001000000000001100000000000,
31'b1010000000000101000000010000000,
31'b0000101000000000000001010000000,
31'b1010000000000001000000010000000,
31'b0000010000000000100000000010000,
31'b0101000000100000010000100000000,
31'b0100000000000000100001001000000,
31'b1010000000001001000000010000000,
31'b0000010000001000100000000010000,
31'b0011010000000100000000100000000,
31'b0001011000000000000000000101000,
31'b0011010000000000000000100000000,
31'b0001000100000000000000010000010,
31'b1000000100000000000001011000000,
31'b1000001000000000000011000100000,
31'b0011010000001000000000100000000,
31'b0001010011000000001000000000000,
31'b1100000000000000000001010100000,
31'b0000101000100000000001010000000,
31'b1010000000100001000000010000000,
31'b0000010000100000100000000010000,
31'b0101000000000000010000100000000,
31'b0101000000000010010000100000000,
31'b0101000000000100010000100000000,
31'b1010000000000000000100000011000,
31'b0100100000001000000011000000000,
31'b0000100000000000000000000011010,
31'b0011010000100000000000100000000,
31'b0001110000000000000001000000001,
31'b0100100000000000000011000000000,
31'b0110000000000000110000000010000,
31'b0001100001000000000000000000010,
31'b1000100000000000000010000001001,
31'b0000000000000000000110000001000,
31'b0000001000000000000000110000010,
31'b0000001000000000010000001100000,
31'b0000010000000000000100001000010,
31'b0000001010100000000001000000000,
31'b0100000010000001000000100001000,
31'b0000100010000000000000000101001,
31'b0001010100010000001000000000000,
31'b0100001000000001000000000010000,
31'b0100001000000011000000000010000,
31'b1100000000000000110010000000000,
31'b0001010100001000001000000000000,
31'b0100001000001001000000000010000,
31'b1010110000000000000000001000000,
31'b0100001100100000010000000000000,
31'b0001010100000000001000000000000,
31'b0000001010001000000001000000000,
31'b0000001010001010000001000000000,
31'b0000100010000000001100001000000,
31'b1100100000000000010000001000000,
31'b0000001010000000000001000000000,
31'b0000001010000010000001000000000,
31'b0000100001000000010010000000000,
31'b1010100010000001000000000000000,
31'b0100001000100001000000000010000,
31'b0000000010000001000100000000010,
31'b1100000000000000000000100010001,
31'b0011000010000000001001000000000,
31'b0100000000000000000010100000010,
31'b0100001000000000000100010001000,
31'b0100001100000000010000000000000,
31'b0100010000000000000000101001000,
31'b0000101000000000001000000000001,
31'b1001000000000000000100000000011,
31'b0000101000000100001000000000001,
31'b0001000010010000000000010000010,
31'b0000101000001000001000000000001,
31'b1100000000000000000100001001000,
31'b0000100000100000010010000000000,
31'b0001000000000000000110000010000,
31'b0110110000000000000010000000000,
31'b1001000000001000000000000100100,
31'b1000000010000000100000100000100,
31'b0001000010000000000000010000010,
31'b1001000000000010000000000100100,
31'b1001000000000000000000000100100,
31'b0001000000100000000001100000000,
31'b0000000000000000110000001000000,
31'b0000101000100000001000000000001,
31'b1100000000000000001000000100001,
31'b0000100000001000010010000000000,
31'b0110100000000000001000000000100,
31'b0000100000000100010010000000000,
31'b0010111000000000000000010000000,
31'b0000100000000000010010000000000,
31'b0010000000000000100001000010000,
31'b1000000000000100010000010100000,
31'b1000000000000000000000101000010,
31'b1000000000000000010000010100000,
31'b1000000000000100000000101000010,
31'b0001000000000100000001100000000,
31'b1001000000100000000000000100100,
31'b0001000000000000000001100000000,
31'b0001000000000010000001100000000,
31'b0000001000101000000001000000000,
31'b0100000000010000000011010000000,
31'b0000100000100000001100001000000,
31'b0001000001010000000000010000010,
31'b0000001000100000000001000000000,
31'b0100000000000001000000100001000,
31'b0000100000000000000000000101001,
31'b1010100000100001000000000000000,
31'b0100001010000001000000000010000,
31'b0100000000000000000011010000000,
31'b1000000001000000100000100000100,
31'b0001000001000000000000010000010,
31'b0000001000110000000001000000000,
31'b0100000000010001000000100001000,
31'b0001100100100000000000000000010,
31'b0001010110000000001000000000000,
31'b0000001000001000000001000000000,
31'b0000001000001010000001000000000,
31'b0000100000000000001100001000000,
31'b1010100000001001000000000000000,
31'b0000001000000000000001000000000,
31'b0000001000000010000001000000000,
31'b0000001000000100000001000000000,
31'b1010100000000001000000000000000,
31'b0000001000011000000001000000000,
31'b0000000000000001000100000000010,
31'b0011000000000010001001000000000,
31'b0011000000000000001001000000000,
31'b0000001000010000000001000000000,
31'b0000001000010010000001000000000,
31'b0001100100000000000000000000010,
31'b1010100000010001000000000000000,
31'b0000101010000000001000000000001,
31'b0001100000000000000000000110001,
31'b1010000100000001000000010000000,
31'b0001000000010000000000010000010,
31'b0000001001100000000001000000000,
31'b0100000100000000100001001000000,
31'b0000100010100000010010000000000,
31'b0001000010000000000110000010000,
31'b1000000000001000000001011000000,
31'b0001000000000100000000010000010,
31'b1000000000000000100000100000100,
31'b0001000000000000000000010000010,
31'b1000000000000000000001011000000,
31'b1001000010000000000000000100100,
31'b1000000000001000100000100000100,
31'b0001000000001000000000010000010,
31'b0000001001001000000001000000000,
31'b0000011000000000000000000000011,
31'b0000100010001000010010000000000,
31'b0001001000000000000001000011000,
31'b0000001001000000000001000000000,
31'b0000010000000001110000000000000,
31'b0000100010000000010010000000000,
31'b1010100001000001000000000000000,
31'b0000000000001000010000000000110,
31'b0000000000000000100001000100000,
31'b1000000010000000010000010100000,
31'b0001000000100000000000010000010,
31'b0000000000000000010000000000110,
31'b0000000000001000100001000100000,
31'b0001000010000000000001100000000,
31'b0001000010000010000001100000000,
31'b0010100000000000000000000000000,
31'b0010100000000010000000000000000,
31'b0010100000000100000000000000000,
31'b1000001000000001000001000000000,
31'b0010100000001000000000000000000,
31'b0010100000001010000000000000000,
31'b1000000000010000000100000000010,
31'b1000001000001001000001000000000,
31'b0010100000010000000000000000000,
31'b0010100000010010000000000000000,
31'b1000000000001000000100000000010,
31'b1000001000010001000001000000000,
31'b1000000000000100000100000000010,
31'b1010001100000000000000001000000,
31'b1000000000000000000100000000010,
31'b1000000000000010000100000000010,
31'b0010100000100000000000000000000,
31'b0000000000000000000001100000001,
31'b1100000000000000000000100001000,
31'b0010000000000001000000000001100,
31'b0010100000101000000000000000000,
31'b0010000101000000000000010000000,
31'b1100000000001000000000100001000,
31'b0010000101000100000000010000000,
31'b0010100000110000000000000000000,
31'b0010000000000000100010001000000,
31'b1100000000010000000000100001000,
31'b0010000000010001000000000001100,
31'b1110000001000000100000000000000,
31'b0010000101010000000000010000000,
31'b1000000000100000000100000000010,
31'b1100001010000000000000000010000,
31'b0010100001000000000000000000000,
31'b0010100001000010000000000000000,
31'b1000010000000000110000000000000,
31'b1000010000000010110000000000000,
31'b0010100001001000000000000000000,
31'b0010000100100000000000010000000,
31'b1000010000001000110000000000000,
31'b0101000100000000001010000000000,
31'b0100010000000000000100000001000,
31'b0110000000000000000000011100000,
31'b1000010000010000110000000000000,
31'b1000010000000000000101000000001,
31'b1110000000100000100000000000000,
31'b0010101000000000100000000100000,
31'b1000000001000000000100000000010,
31'b1000001000000000100000000000101,
31'b0010100001100000000000000000000,
31'b0010000100001000000000010000000,
31'b1100000001000000000000100001000,
31'b0010000100001100000000010000000,
31'b0000010000000000000000100000010,
31'b0010000100000000000000010000000,
31'b0010000000000000010100000001000,
31'b0010000100000100000000010000000,
31'b1110000000001000100000000000000,
31'b0010000100011000000000010000000,
31'b0001001100000000001000010000000,
31'b0000000100000000000010000000101,
31'b1110000000000000100000000000000,
31'b0010000100010000000000010000000,
31'b1110000000000100100000000000000,
31'b0010000100010100000000010000000,
31'b0010100010000000000000000000000,
31'b0010100010000010000000000000000,
31'b1000000000000000000010010010000,
31'b1000001010000001000001000000000,
31'b0000000000000000000000010000011,
31'b0000100001000000001000100000000,
31'b0000100000010000000000000110000,
31'b0100000001000000000000011010000,
31'b0010100010010000000000000000000,
31'b0010100010010010000000000000000,
31'b0010000000000000000010000000110,
31'b0100000100000000100010000010000,
31'b0000100000000100000000000110000,
31'b0100000000000100011000000000010,
31'b0000100000000000000000000110000,
31'b0100000000000000011000000000010,
31'b0010100010100000000000000000000,
31'b0010010000000000001000000000010,
31'b1100000010000000000000100001000,
31'b0010010000000100001000000000010,
31'b0000110100000000000001000000000,
31'b0010010000001000001000000000010,
31'b0001011000010000000000000000010,
31'b1100001000010000000000000010000,
31'b0010100010110000000000000000000,
31'b1100000000000000101000100000000,
31'b0010110000000001000000001000000,
31'b1100001000001000000000000010000,
31'b0001011000000100000000000000010,
31'b1100001000000100000000000010000,
31'b0001011000000000000000000000010,
31'b1100001000000000000000000010000,
31'b0010100011000000000000000000000,
31'b0000010000000000000001010000000,
31'b1000010010000000110000000000000,
31'b0000101000000000100000000010000,
31'b0000100000000010001000100000000,
31'b0000100000000000001000100000000,
31'b0100000000000010000000011010000,
31'b0100000000000000000000011010000,
31'b0111000000000000000001000000100,
31'b0001100000000000000000000101000,
31'b0011101000000000000000100000000,
31'b0001100000000100000000000101000,
31'b0000100001000100000000000110000,
31'b0000100000010000001000100000000,
31'b0000100001000000000000000110000,
31'b0100000001000000011000000000010,
31'b0010100011100000000000000000000,
31'b0000100100000000000000000000011,
31'b1100000000000000100000000110000,
31'b0001010000000000100000000100010,
31'b0010000000000000001001000000001,
31'b0010000110000000000000010000000,
31'b0010000010000000010100000001000,
31'b1110000000000000001000000001000,
31'b1101001000000000000000000001000,
31'b0001100000100000000000000101000,
31'b0001000000000001000000000100100,
31'b0001001000000000000001000000001,
31'b1110000010000000100000000000000,
31'b0010000110010000000000010000000,
31'b0001011001000000000000000000010,
31'b1100001001000000000000000010000,
31'b0010100100000000000000000000000,
31'b0010100100000010000000000000000,
31'b1001000000000000001000001000000,
31'b1001000000000010001000001000000,
31'b0010100100001000000000000000000,
31'b0000000000000000001001000000010,
31'b1001000000001000001000001000000,
31'b0011000000000001000100000000000,
31'b0010100100010000000000000000000,
31'b1010001000001000000000001000000,
31'b1001000000010000001000001000000,
31'b0100010001000000010000010000000,
31'b1010001000000010000000001000000,
31'b1010001000000000000000001000000,
31'b1000000100000000000100000000010,
31'b1010001000000100000000001000000,
31'b0010100100100000000000000000000,
31'b0010000001001000000000010000000,
31'b1100000100000000000000100001000,
31'b0010000100000001000000000001100,
31'b0010000001000010000000010000000,
31'b0010000001000000000000010000000,
31'b0010100000000001010000000010000,
31'b0010000001000100000000010000000,
31'b0010100100110000000000000000000,
31'b0010000100000000100010001000000,
31'b1001000000000000000000000001110,
31'b0000000001000000000010000000101,
31'b0110100000000000000000001100000,
31'b0010000001010000000000010000000,
31'b1100000000000000000000001000101,
31'b0010000001010100000000010000000,
31'b0000010000000000001000000000001,
31'b0010000000101000000000010000000,
31'b0011000000000000010000000000100,
31'b0101000000001000001010000000000,
31'b0010000000100010000000010000000,
31'b0010000000100000000000010000000,
31'b0101000000000010001010000000000,
31'b0101000000000000001010000000000,
31'b0110001000000000000010000000000,
31'b0110001000000010000010000000000,
31'b0110001000000100000010000000000,
31'b0100010000000000010000010000000,
31'b0110001000001000000010000000000,
31'b0010000000110000000000010000000,
31'b1000000101000000000100000000010,
31'b0101000000010000001010000000000,
31'b0010000000001010000000010000000,
31'b0010000000001000000000010000000,
31'b0011000000100000010000000000100,
31'b0010000000001100000000010000000,
31'b0010000000000010000000010000000,
31'b0010000000000000000000010000000,
31'b0010000000000110000000010000000,
31'b0010000000000100000000010000000,
31'b0110001000100000000010000000000,
31'b0010000000011000000000010000000,
31'b0001001000000000001000010000000,
31'b0000000000000000000010000000101,
31'b0101010000000000000000000000100,
31'b0010000000010000000000010000000,
31'b0110000000000000011000000000001,
31'b0010000000010100000000010000000,
31'b0010100110000000000000000000000,
31'b0010100110000010000000000000000,
31'b1001000010000000001000001000000,
31'b1001000000000001000010000000100,
31'b0000110000100000000001000000000,
31'b0010010000000000000000100000001,
31'b0000110000100100000001000000000,
31'b0011000010000001000100000000000,
31'b0010100110010000000000000000000,
31'b1100001000000001010000000000000,
31'b0110100000000000010001000000000,
31'b0100000000000000100010000010000,
31'b0001010000000000100000000010001,
31'b1100000000000000100000000000011,
31'b0000100100000000000000000110000,
31'b0100000100000000011000000000010,
31'b0000000000000000001000110000000,
31'b0000100001000000000000000000011,
31'b0100100000000000000000001010000,
31'b0100100000000010000000001010000,
31'b0000110000000000000001000000000,
31'b0010000011000000000000010000000,
31'b0000110000000100000001000000000,
31'b1010011000000001000000000000000,
31'b0000100000000001010000000100000,
31'b0100000000000100010000100000001,
31'b0100100000010000000000001010000,
31'b0100000000000000010000100000001,
31'b0001000000000000000000010101000,
31'b0011010000000000000100001000000,
31'b0001011100000000000000000000010,
31'b1100001100000000000000000010000,
31'b0010000000000000000001100000010,
31'b0000100000100000000000000000011,
31'b0011000010000000010000000000100,
31'b0000101100000000100000000010000,
31'b0010000010100010000000010000000,
31'b0010000010100000000000010000000,
31'b1001000000000000010110000000000,
31'b1011000000000000000000101000000,
31'b1100010000000000100001000000000,
31'b0001100100000000000000000101000,
31'b1000010000000000001100010000000,
31'b0000010000000000100000000001001,
31'b1100001000000000000100000000100,
31'b0010001000000001000100100000000,
31'b1000000000000000100000001010000,
31'b1010000000100000000100000000001,
31'b0000100000000010000000000000011,
31'b0000100000000000000000000000011,
31'b0100100001000000000000001010000,
31'b0000100000000100000000000000011,
31'b0010000010000010000000010000000,
31'b0010000010000000000000010000000,
31'b1010000000000000110001000000000,
31'b1000100000000000000010000010000,
31'b0000100001000001010000000100000,
31'b0000100000010000000000000000011,
31'b0000000000000010000000010110000,
31'b0000000000000000000000010110000,
31'b0110000000000000000101000001000,
31'b0010000010010000000000010000000,
31'b1010000000000010000100000000001,
31'b1010000000000000000100000000001,
31'b0010101000000000000000000000000,
31'b1000000000000101000001000000000,
31'b1000000000000011000001000000000,
31'b1000000000000001000001000000000,
31'b0010101000001000000000000000000,
31'b1010000100010000000000001000000,
31'b1000001000010000000100000000010,
31'b1000000000001001000001000000000,
31'b0010101000010000000000000000000,
31'b1010000100001000000000001000000,
31'b1000001000001000000100000000010,
31'b1000000000010001000001000000000,
31'b1010000100000010000000001000000,
31'b1010000100000000000000001000000,
31'b1000001000000000000100000000010,
31'b0001100000000000001000000000000,
31'b0010101000100000000000000000000,
31'b1110000000000000000000000100000,
31'b1100001000000000000000100001000,
31'b1000000000100001000001000000000,
31'b0010101000101000000000000000000,
31'b1110000000001000000000000100000,
31'b0001010010010000000000000000010,
31'b1100000010010000000000000010000,
31'b0010101000110000000000000000000,
31'b1110000000010000000000000100000,
31'b0001010010001000000000000000010,
31'b1100000010001000000000000010000,
31'b0001010010000100000000000000010,
31'b1100000010000100000000000010000,
31'b0001010010000000000000000000010,
31'b1100000010000000000000000010000,
31'b0010101001000000000000000000000,
31'b1010000000000000100010010000000,
31'b1000011000000000110000000000000,
31'b1000000001000001000001000000000,
31'b0010101001001000000000000000000,
31'b0010100000010000100000000100000,
31'b1000010000000001000000000000011,
31'b1000000001001001000001000000000,
31'b0110000100000000000010000000000,
31'b0110000100000010000010000000000,
31'b0110000100000100000010000000000,
31'b1000000001010001000001000000000,
31'b0110000100001000000010000000000,
31'b0010100000000000100000000100000,
31'b1000001001000000000100000000010,
31'b1000000000000000100000000000101,
31'b0010101001100000000000000000000,
31'b1110000001000000000000000100000,
31'b0001000100010000001000010000000,
31'b1101000000000000101000000000000,
31'b0010000000000000000010001100000,
31'b0010001100000000000000010000000,
31'b0000010100000000010010000000000,
31'b0010010000000000000000000101010,
31'b1101000010000000000000000001000,
31'b0001000010000100000001000000001,
31'b0001000100000000001000010000000,
31'b0001000010000000000001000000001,
31'b1110001000000000100000000000000,
31'b0010100000100000100000000100000,
31'b0001010011000000000000000000010,
31'b1100000011000000000000000010000,
31'b0010101010000000000000000000000,
31'b1010010000000000010000000010000,
31'b1000001000000000000010010010000,
31'b1000000010000001000001000000000,
31'b0001100000000000100000000001000,
31'b0001100000000010100000000001000,
31'b0001100000000100100000000001000,
31'b1100000000110000000000000010000,
31'b0010101010010000000000000000000,
31'b1100000100000001010000000000000,
31'b0011100001000000000000100000000,
31'b1100000000101000000000000010000,
31'b0001100000010000100000000001000,
31'b1100000000100100000000000010000,
31'b0001010000100000000000000000010,
31'b1100000000100000000000000010000,
31'b0010101010100000000000000000000,
31'b1110000010000000000000000100000,
31'b0001010000011000000000000000010,
31'b1100000000011000000000000010000,
31'b0001100000100000100000000001000,
31'b1100000000010100000000000010000,
31'b0001010000010000000000000000010,
31'b1100000000010000000000000010000,
31'b1101000001000000000000000001000,
31'b1000010000000000000001001000000,
31'b0001010000001000000000000000010,
31'b1100000000001000000000000010000,
31'b0001010000000100000000000000010,
31'b1100000000000100000000000010000,
31'b0001010000000000000000000000010,
31'b1100000000000000000000000010000,
31'b0010101011000000000000000000000,
31'b0000100000000100100000000010000,
31'b0010000000000000010011000000000,
31'b0000100000000000100000000010000,
31'b1001000000000000000100100000010,
31'b0000101000000000001000100000000,
31'b0100000100000000000010000110000,
31'b0100000000000000001001000000100,
31'b1101000000100000000000000001000,
31'b0001101000000000000000000101000,
31'b0011100000000000000000100000000,
31'b0001000000100000000001000000001,
31'b1100000100000000000100000000100,
31'b0010100010000000100000000100000,
31'b0011100000001000000000100000000,
31'b1100000001100000000000000010000,
31'b1101000000010000000000000001000,
31'b0001000100000000100000010001000,
31'b0001000000000000110100000000000,
31'b0001000000010000000001000000001,
31'b1100000000000000001000100100000,
31'b0010001110000000000000010000000,
31'b0001010001010000000000000000010,
31'b1100000001010000000000000010000,
31'b1101000000000000000000000001000,
31'b0001000000000100000001000000001,
31'b0000000000000000000010001010000,
31'b0001000000000000000001000000001,
31'b1000000000000000000000001000011,
31'b1100000001000100000000000010000,
31'b0001010001000000000000000000010,
31'b1100000001000000000000000010000,
31'b0010101100000000000000000000000,
31'b1010000000011000000000001000000,
31'b1001001000000000001000001000000,
31'b1000000100000001000001000000000,
31'b1010000000010010000000001000000,
31'b1010000000010000000000001000000,
31'b0100000001000000000000010000101,
31'b1010000000010100000000001000000,
31'b0000000000000001001100000000000,
31'b1010000000001000000000001000000,
31'b0011000000000000000001000000010,
31'b1010000000001100000000001000000,
31'b1010000000000010000000001000000,
31'b1010000000000000000000001000000,
31'b1010000000000110000000001000000,
31'b1010000000000100000000001000000,
31'b0010101100100000000000000000000,
31'b1110000100000000000000000100000,
31'b0001000001010000001000010000000,
31'b1100010000000000010000001000000,
31'b1010100000000000100010000000000,
31'b1000000000000000010001000010000,
31'b0000010001000000010010000000000,
31'b1010010010000001000000000000000,
31'b0010000000000000100000010100000,
31'b1010000000101000000000001000000,
31'b0001000001000000001000010000000,
31'b0001100000000000000000100000011,
31'b1010000000100010000000001000000,
31'b1010000000100000000000001000000,
31'b0001010110000000000000000000010,
31'b1100000110000000000000000010000,
31'b0110000000010000000010000000000,
31'b0110000000010010000010000000000,
31'b0110000000010100000010000000000,
31'b1000000101000001000001000000000,
31'b0110000000011000000010000000000,
31'b0010001000100000000000010000000,
31'b0100000000000000000000010000101,
31'b0101001000000000001010000000000,
31'b0110000000000000000010000000000,
31'b0110000000000010000010000000000,
31'b0110000000000100000010000000000,
31'b0110000000000110000010000000000,
31'b0110000000001000000010000000000,
31'b0000000000000000011000000000100,
31'b0110000000001100000010000000000,
31'b0011010000000000000000000000001,
31'b0110000000110000000010000000000,
31'b0101000000000000010000000000001,
31'b0001000000010000001000010000000,
31'b0110010000000000001000000000100,
31'b0010001000000010000000010000000,
31'b0010001000000000000000010000000,
31'b0000010000000000010010000000000,
31'b0010001000000100000000010000000,
31'b0110000000100000000010000000000,
31'b0110000000100010000010000000000,
31'b0001000000000000001000010000000,
31'b0001000000000010001000010000000,
31'b0110000000101000000010000000000,
31'b0010001000010000000000010000000,
31'b0001000000001000001000010000000,
31'b0011010000100000000000000000001,
31'b0010101110000000000000000000000,
31'b1100000000010001010000000000000,
31'b1000000000000010000000001110000,
31'b1000000000000000000000001110000,
31'b0001100100000000100000000001000,
31'b1100010000000000000001000100000,
31'b0000010000000000000000000101001,
31'b1010010000100001000000000000000,
31'b0010000000000000010000100000100,
31'b1100000000000001010000000000000,
31'b0011000010000000000001000000010,
31'b1100000000000101010000000000000,
31'b1100000001000000000100000000100,
31'b1010000010000000000000001000000,
31'b0001100000000000000001010000001,
31'b1100000100100000000000000010000,
31'b0000100000000000100100000000100,
31'b0001000001000000100000010001000,
31'b0000010000000000001100001000000,
31'b1010010000001001000000000000000,
31'b0000111000000000000001000000000,
31'b1010010000000101000000000000000,
31'b0000000000000000100000010010000,
31'b1010010000000001000000000000000,
31'b0010000010000000100000010100000,
31'b1100000000100001010000000000000,
31'b0001010100001000000000000000010,
31'b1100000100001000000000000010000,
31'b0001010100000100000000000000010,
31'b1100000100000100000000000010000,
31'b0001010100000000000000000000010,
31'b1100000100000000000000000010000,
31'b1100000000000000000000000100011,
31'b0001010000000000000000000110001,
31'b0110100000000000000000000000110,
31'b0000100100000000100000000010000,
31'b1100000000010000000100000000100,
31'b0010001010100000000000010000000,
31'b0100000000000000000010000110000,
31'b0100000100000000001001000000100,
31'b1000000000000000001000101000000,
31'b1100000001000001010000000000000,
31'b1100100000000000000000010010000,
31'b0001110000000000000000010000010,
31'b1100000000000000000100000000100,
31'b0010000000000001000100100000000,
31'b1100000000000100000100000000100,
31'b0011010010000000000000000000001,
31'b1001000000000000001100000000001,
31'b0001000000000000100000010001000,
31'b0001000100000000110100000000000,
31'b0001000100010000000001000000001,
31'b0010001010000010000000010000000,
31'b0010001010000000000000010000000,
31'b0000010010000000010010000000000,
31'b1010010001000001000000000000000,
31'b1101000100000000000000000001000,
31'b0001000100000100000001000000001,
31'b0001000010000000001000010000000,
31'b0001000100000000000001000000001,
31'b1100000000100000000100000000100,
31'b0010001010010000000000010000000,
31'b0001010101000000000000000000010,
31'b1100000101000000000000000010000,
31'b0010110000000000000000000000000,
31'b0010110000000010000000000000000,
31'b1000000001000000110000000000000,
31'b1000011000000001000001000000000,
31'b0010110000001000000000000000000,
31'b0010110000001010000000000000000,
31'b1000010000010000000100000000010,
31'b1000001000010000010000000100000,
31'b0100000001000000000100000001000,
31'b0101100000000000000000010000100,
31'b1000010000001000000100000000010,
31'b1000001000001000010000000100000,
31'b1010000000000000010000100001000,
31'b1000001000000100010000000100000,
31'b1000010000000000000100000000010,
31'b1000001000000000010000000100000,
31'b0010110000100000000000000000000,
31'b0010000010000000001000000000010,
31'b1100010000000000000000100001000,
31'b0010010000000001000000000001100,
31'b0000000001000000000000100000010,
31'b0000100000000000001000010000001,
31'b0100100000010000010000000000000,
31'b0100100000010010010000000000000,
31'b0100100000001100010000000000000,
31'b1000001010000000000001001000000,
31'b0100100000001000010000000000000,
31'b0100100000001010010000000000000,
31'b0100100000000100010000000000000,
31'b0100100000000110010000000000000,
31'b0100100000000000010000000000000,
31'b0100100000000010010000000000000,
31'b0000000100000000001000000000001,
31'b0000000010000000000001010000000,
31'b1000000000000000110000000000000,
31'b1000000000000010110000000000000,
31'b0000000000100000000000100000010,
31'b0000000010001000000001010000000,
31'b1000000000001000110000000000000,
31'b1000000000001010110000000000000,
31'b0100000000000000000100000001000,
31'b0100000000000010000100000001000,
31'b1000000000010000110000000000000,
31'b1000000000000000000101000000001,
31'b0100000000001000000100000001000,
31'b0100000000100001000000010010000,
31'b1000010001000000000100000000010,
31'b1000001001000000010000000100000,
31'b0000000000001000000000100000010,
31'b0000000010100000000001010000000,
31'b1000000000100000110000000000000,
31'b1001000000000000000001101000000,
31'b0000000000000000000000100000010,
31'b0000000000000010000000100000010,
31'b0000000000000100000000100000010,
31'b0000000000000110000000100000010,
31'b0100000000100000000100000001000,
31'b0100000000100010000100000001000,
31'b1010100000000000000100100000000,
31'b1000100000000000010010001000000,
31'b0000000000010000000000100000010,
31'b0100000000000001000000010010000,
31'b0100100001000000010000000000000,
31'b0100100001000010010000000000000,
31'b0010110010000000000000000000000,
31'b0000000001000000000001010000000,
31'b1000010000000000000010010010000,
31'b0010000000000001100010000000000,
31'b0000100100100000000001000000000,
31'b0010000100000000000000100000001,
31'b0001001000110000000000000000010,
31'b0010000100000100000000100000001,
31'b0100100000000000000001001100000,
31'b0010000000000000000000001001100,
31'b0010100000100001000000001000000,
31'b0010000000010001100010000000000,
31'b0001001000100100000000000000010,
31'b0010000100010000000000100000001,
31'b0001001000100000000000000000010,
31'b1000100000100000001100000000000,
31'b0010000000000010001000000000010,
31'b0010000000000000001000000000010,
31'b0010100000010001000000001000000,
31'b0010000000000100001000000000010,
31'b0000100100000000000001000000000,
31'b0010000000001000001000000000010,
31'b0001001000010000000000000000010,
31'b1010001100000001000000000000000,
31'b1001000100000001001000000000000,
31'b1000001000000000000001001000000,
31'b0010100000000001000000001000000,
31'b1000100000001000001100000000000,
31'b0001001000000100000000000000010,
31'b1000100000000100001100000000000,
31'b0001001000000000000000000000010,
31'b1000100000000000001100000000000,
31'b0000000000000010000001010000000,
31'b0000000000000000000001010000000,
31'b1000000010000000110000000000000,
31'b0000000000000100000001010000000,
31'b0000000010100000000000100000010,
31'b0000000000001000000001010000000,
31'b1001000000000000000000011000010,
31'b0000000000001100000001010000000,
31'b0100000010000000000100000001000,
31'b0000000000010000000001010000000,
31'b1000000100000000001100010000000,
31'b0000000100000000100000000001001,
31'b0100001000100000000011000000000,
31'b0000000000011000000001010000000,
31'b0011000000000000000000001010100,
31'b0010000100000001000000011000000,
31'b0000000010001000000000100000010,
31'b0000000000100000000001010000000,
31'b1000000010100000110000000000000,
31'b0001000000000000100000000100010,
31'b0000000010000000000000100000010,
31'b0000000010000010000000100000010,
31'b0001000000000000010001000000100,
31'b0001000000001000100000000100010,
31'b0100001000001000000011000000000,
31'b0000001000000000000000000011010,
31'b0010100001000001000000001000000,
31'b0001011000000000000001000000001,
31'b0100001000000000000011000000000,
31'b0100001000000010000011000000000,
31'b0001001001000000000000000000010,
31'b1000100001000000001100000000000,
31'b0000000001000000001000000000001,
31'b0000100000000000000000110000010,
31'b0000100000000000010000001100000,
31'b0100000001010000010000010000000,
31'b0000100010100000000001000000000,
31'b0010000010000000000000100000001,
31'b0000100010100100000001000000000,
31'b0011010000000001000100000000000,
31'b0100100000000001000000000010000,
31'b0100100000000011000000000010000,
31'b0100100000000101000000000010000,
31'b0100000001000000010000010000000,
31'b0101000001100000000000000000100,
31'b1010011000000000000000001000000,
31'b1000010100000000000100000000010,
31'b1010000000000000000100110000000,
31'b0000100010001000000001000000000,
31'b0010010001001000000000010000000,
31'b0000100010001100000001000000000,
31'b1100001000000000010000001000000,
31'b0000100010000000000001000000000,
31'b0010010001000000000000010000000,
31'b0000100010000100000001000000000,
31'b1010001010000001000000000000000,
31'b1001000010000001001000000000000,
31'b1001000000000000000010001000100,
31'b0100100100001000010000000000000,
31'b0100000000000000000000000011100,
31'b0101000001000000000000000000100,
31'b0101000001000010000000000000100,
31'b0100100100000000010000000000000,
31'b0100100100000010010000000000000,
31'b0000000000000000001000000000001,
31'b0000000000000010001000000000001,
31'b0000000000000100001000000000001,
31'b0100000000010000010000010000000,
31'b0000000000001000001000000000001,
31'b0010010000100000000000010000000,
31'b0000001000100000010010000000000,
31'b0101010000000000001010000000000,
31'b0000000000010000001000000000001,
31'b0100000000000100010000010000000,
31'b0100000000000010010000010000000,
31'b0100000000000000010000010000000,
31'b0101000000100000000000000000100,
31'b0101000000100010000000000000100,
31'b0101000000100100000000000000100,
31'b0100000000001000010000010000000,
31'b0000000000100000001000000000001,
31'b0010010000001000000000010000000,
31'b0000001000001000010010000000000,
31'b0110001000000000001000000000100,
31'b0000000100000000000000100000010,
31'b0010010000000000000000010000000,
31'b0000001000000000010010000000000,
31'b0010010000000100000000010000000,
31'b0101000000001000000000000000100,
31'b0101000000001010000000000000100,
31'b0101000000001100000000000000100,
31'b0100000000100000010000010000000,
31'b0101000000000000000000000000100,
31'b0101000000000010000000000000100,
31'b0101000000000100000000000000100,
31'b0101000000000110000000000000100,
31'b0000100000101000000001000000000,
31'b0010000000001000000000100000001,
31'b0000100010000000010000001100000,
31'b0010000100000001100010000000000,
31'b0000100000100000000001000000000,
31'b0010000000000000000000100000001,
31'b0000100000100100000001000000000,
31'b0010000000000100000000100000001,
31'b1100000001000000100001000000000,
31'b0010000100000000000000001001100,
31'b1001000000000000100010000000010,
31'b0000000001000000100000000001001,
31'b0001000000000000100000000010001,
31'b0010000000010000000000100000001,
31'b0001001100100000000000000000010,
31'b0010000001000001000000011000000,
31'b0000100000001000000001000000000,
31'b0010000100000000001000000000010,
31'b0000100000001100000001000000000,
31'b1010001000001001000000000000000,
31'b0000100000000000000001000000000,
31'b0000100000000010000001000000000,
31'b0000100000000100000001000000000,
31'b1010001000000001000000000000000,
31'b1001000000000001001000000000000,
31'b1001000000000011001000000000000,
31'b1010000000000000000101000000010,
31'b0100010000000000010000100000001,
31'b0000100000010000000001000000000,
31'b0011000000000000000100001000000,
31'b0001001100000000000000000000010,
31'b1010001000010001000000000000000,
31'b0000000010000000001000000000001,
31'b0000000100000000000001010000000,
31'b0000000010000100001000000000001,
31'b0000000100000100000001010000000,
31'b0000100001100000000001000000000,
31'b0010000001000000000000100000001,
31'b0000100001100100000001000000000,
31'b0010000001000100000000100000001,
31'b1100000000000000100001000000000,
31'b0000000100010000000001010000000,
31'b1000000000000000001100010000000,
31'b0000000000000000100000000001001,
31'b1100000000001000100001000000000,
31'b0010000001010000000000100000001,
31'b1000010000000000100000001010000,
31'b0010000000000001000000011000000,
31'b0000100001001000000001000000000,
31'b0000110000000000000000000000011,
31'b0000100001001100000001000000000,
31'b0001100000000000000001000011000,
31'b0000100001000000000001000000000,
31'b0010010010000000000000010000000,
31'b0000100001000100000001000000000,
31'b1010001001000001000000000000000,
31'b1100000000100000100001000000000,
31'b0000110000010000000000000000011,
31'b1010000000000001100000000100000,
31'b0000010000000000000000010110000,
31'b0101000010000000000000000000100,
31'b0101000010000010000000000000100,
31'b0101000010000100000000000000100,
31'b1010010000000000000100000000001,
31'b0010111000000000000000000000000,
31'b1010000010000000010000000010000,
31'b1000010000000011000001000000000,
31'b1000010000000001000001000000000,
31'b0010111000001000000000000000000,
31'b1100000000000001000000001010000,
31'b1000000001000001000000000000011,
31'b1000000000010000010000000100000,
31'b0100100000000000001010000000001,
31'b1000000010100000000001001000000,
31'b1000000000001010010000000100000,
31'b1000000000001000010000000100000,
31'b1000000000000110010000000100000,
31'b1000000000000100010000000100000,
31'b1000000000000010010000000100000,
31'b1000000000000000010000000100000,
31'b0011000000000000000000000110010,
31'b1110010000000000000000000100000,
31'b0001000010011000000000000000010,
31'b1100000100000000010000001000000,
31'b0001100000000000000010000000100,
31'b0001100000000010000010000000100,
31'b0001000010010000000000000000010,
31'b1010000110000001000000000000000,
31'b1001000000000000000000010100100,
31'b1000000010000000000001001000000,
31'b0001000010001000000000000000010,
31'b1000000010000100000001001000000,
31'b0001000010000100000000000000010,
31'b1000000010001000000001001000000,
31'b0001000010000000000000000000010,
31'b1000000000100000010000000100000,
31'b0000000000000001000010000010000,
31'b0000001010000000000001010000000,
31'b1000001000000000110000000000000,
31'b1000010001000001000001000000000,
31'b0000001000100000000000100000010,
31'b0100000010000000000100100010000,
31'b1000000000000001000000000000011,
31'b1000000001010000010000000100000,
31'b0100001000000000000100000001000,
31'b0100001000000010000100000001000,
31'b1000001000010000110000000000000,
31'b1000001000000000000101000000001,
31'b0100001000001000000100000001000,
31'b1000100000000000001000001000001,
31'b1000000001000010010000000100000,
31'b1000000001000000010000000100000,
31'b0000001000001000000000100000010,
31'b0000001010100000000001010000000,
31'b0000000100001000010010000000000,
31'b0110000100000000001000000000100,
31'b0000001000000000000000100000010,
31'b0000001000000010000000100000010,
31'b0000000100000000010010000000000,
31'b0010000000000000000000000101010,
31'b0100001000100000000100000001000,
31'b0000000010000000000000000011010,
31'b0001010100000000001000010000000,
31'b0011000000000000001000100000010,
31'b0100000010000000000011000000000,
31'b0100001000000001000000010010000,
31'b0001000011000000000000000000010,
31'b1000000010000000000010000001001,
31'b1010000000000010010000000010000,
31'b1010000000000000010000000010000,
31'b0101000000000000000100100001000,
31'b1010000000000100010000000010000,
31'b0001110000000000100000000001000,
31'b1100000100000000000001000100000,
31'b0001000000110000000000000000010,
31'b1010000100100001000000000000000,
31'b1001000000000000110000100000000,
31'b1000000000100000000001001000000,
31'b0001000000101000000000000000010,
31'b1000000010001000010000000100000,
31'b0001000000100100000000000000010,
31'b1000000010000100010000000100000,
31'b0001000000100000000000000000010,
31'b1000000010000000010000000100000,
31'b1011100000000000000100000000000,
31'b1000000000010000000001001000000,
31'b0001000000011000000000000000010,
31'b1010000100001001000000000000000,
31'b0001000000010100000000000000010,
31'b1010000100000101000000000000000,
31'b0001000000010000000000000000010,
31'b1010000100000001000000000000000,
31'b1000000000000010000001001000000,
31'b1000000000000000000001001000000,
31'b0001000000001000000000000000010,
31'b1000000000000100000001001000000,
31'b0001000000000100000000000000010,
31'b1000000000001000000001001000000,
31'b0001000000000000000000000000010,
31'b0001000000000010000000000000010,
31'b0000001000000010000001010000000,
31'b0000001000000000000001010000000,
31'b1010100000000001000000010000000,
31'b0000110000000000100000000010000,
31'b0100000000110000000011000000000,
31'b0100000000000000000100100010000,
31'b1011000000000000010000000001000,
31'b0100010000000000001001000000100,
31'b0100001010000000000100000001000,
31'b0000001000010000000001010000000,
31'b0011110000000000000000100000000,
31'b0001100100000000000000010000010,
31'b0100000000100000000011000000000,
31'b0100000000100010000011000000000,
31'b0010000000000001000010000100000,
31'b1000000011000000010000000100000,
31'b0100000000011000000011000000000,
31'b0000001000100000000001010000000,
31'b0001010000000000110100000000000,
31'b0001010000010000000001000000001,
31'b0100000000010000000011000000000,
31'b0100000000100000000100100010000,
31'b0001000001010000000000000000010,
31'b1010000101000001000000000000000,
31'b0100000000001000000011000000000,
31'b0000000000000000000000000011010,
31'b0001000001001000000000000000010,
31'b0001010000000000000001000000001,
31'b0100000000000000000011000000000,
31'b0100000000000010000011000000000,
31'b0001000001000000000000000000010,
31'b1000000000000000000010000001001,
31'b0000100000000000000110000001000,
31'b0001000001000000000010010000100,
31'b0000101000000000010000001100000,
31'b1100000000100000010000001000000,
31'b0000101010100000000001000000000,
31'b1100000010000000000001000100000,
31'b0000000010000000000000000101001,
31'b1010000010100001000000000000000,
31'b0010000000000000000000000011001,
31'b1010010000001000000000001000000,
31'b0011010000000000000001000000010,
31'b1110000000000000000001000010000,
31'b1010010000000010000000001000000,
31'b1010010000000000000000001000000,
31'b1010000000000000000010000001010,
31'b1000000100000000010000000100000,
31'b0000101010001000000001000000000,
31'b1100000000000100010000001000000,
31'b0000000010000000001100001000000,
31'b1100000000000000010000001000000,
31'b0000101010000000000001000000000,
31'b1010000010000101000000000000000,
31'b0000000001000000010010000000000,
31'b1010000010000001000000000000000,
31'b1000000000000011000000000110000,
31'b1000000000000001000000000110000,
31'b0001010001000000001000010000000,
31'b1100000000010000010000001000000,
31'b0101001001000000000000000000100,
31'b1010010000100000000000001000000,
31'b0001000110000000000000000000010,
31'b1010000010010001000000000000000,
31'b0000001000000000001000000000001,
31'b0001000000000000000010010000100,
31'b0000001000000100001000000000001,
31'b0110000000100000001000000000100,
31'b0000001000001000001000000000001,
31'b0011000000010100000000000000001,
31'b0000000000100000010010000000000,
31'b0011000000010000000000000000001,
31'b0110010000000000000010000000000,
31'b0110010000000010000010000000000,
31'b0110010000000100000010000000000,
31'b0100001000000000010000010000000,
31'b0110010000001000000010000000000,
31'b0011000000000100000000000000001,
31'b0011000000000010000000000000001,
31'b0011000000000000000000000000001,
31'b0000001000100000001000000000001,
31'b0110000000000100001000000000100,
31'b0000000000001000010010000000000,
31'b0110000000000000001000000000100,
31'b0000000000000100010010000000000,
31'b0010011000000000000000010000000,
31'b0000000000000000010010000000000,
31'b0000000000000010010010000000000,
31'b0110010000100000000010000000000,
31'b1000100000000000000000101000010,
31'b0001010000000000001000010000000,
31'b0110000000010000001000000000100,
31'b0101001000000000000000000000100,
31'b0101001000000010000000000000100,
31'b0000000000010000010010000000000,
31'b0011000000100000000000000000001,
31'b0000101000101000000001000000000,
31'b1100000000001000000001000100000,
31'b0000000000100000001100001000000,
31'b1010000000101001000000000000000,
31'b0000101000100000000001000000000,
31'b1100000000000000000001000100000,
31'b0000000000000000000000000101001,
31'b1010000000100001000000000000000,
31'b0010010000000000010000100000100,
31'b1100010000000001010000000000000,
31'b0001000000000000001000100000001,
31'b0001100001000000000000010000010,
31'b0001001000000000100000000010001,
31'b1100000000010000000001000100000,
31'b0001000100100000000000000000010,
31'b1010000000110001000000000000000,
31'b0000101000001000000001000000000,
31'b1010000000001101000000000000000,
31'b0000000000000000001100001000000,
31'b1010000000001001000000000000000,
31'b0000101000000000000001000000000,
31'b1010000000000101000000000000000,
31'b0100000000000000000000100000100,
31'b1010000000000001000000000000000,
31'b1001001000000001001000000000000,
31'b1000000100000000000001001000000,
31'b0001000100001000000000000000010,
31'b1010000000011001000000000000000,
31'b0001000100000100000000000000010,
31'b1010000000010101000000000000000,
31'b0001000100000000000000000000010,
31'b1010000000010001000000000000000,
31'b0000001010000000001000000000001,
31'b0001000000000000000000000110001,
31'b0000001010000100001000000000001,
31'b0001100000010000000000010000010,
31'b0000101001100000000001000000000,
31'b1100000001000000000001000100000,
31'b0000000010100000010010000000000,
31'b1010000001100001000000000000000,
31'b1100001000000000100001000000000,
31'b0001100000000100000000010000010,
31'b1000100000000000100000100000100,
31'b0001100000000000000000010000010,
31'b1100010000000000000100000000100,
31'b0011000010000100000000000000001,
31'b0011000010000010000000000000001,
31'b0011000010000000000000000000001,
31'b0000101001001000000001000000000,
31'b0001010000000000100000010001000,
31'b0000000010001000010010000000000,
31'b1010000001001001000000000000000,
31'b0000101001000000000001000000000,
31'b1010000001000101000000000000000,
31'b0000000010000000010010000000000,
31'b1010000001000001000000000000000,
31'b0110000000000000100000000001100,
31'b0000100000000000100001000100000,
31'b0001010010000000001000010000000,
31'b0001100000100000000000010000010,
31'b0100000100000000000011000000000,
31'b0100000100000010000011000000000,
31'b0001000101000000000000000000010,
31'b1010000001010001000000000000000,
31'b0011000000000000000000000000000,
31'b0011000000000010000000000000000,
31'b0011000000000100000000000000000,
31'b0011000000000110000000000000000,
31'b0011000000001000000000000000000,
31'b0011000000001010000000000000000,
31'b0011000000001100000000000000000,
31'b0000001000010000001000000000000,
31'b0011000000010000000000000000000,
31'b0000000000000000100000100010000,
31'b0011000000010100000000000000000,
31'b0000001000001000001000000000000,
31'b0011000000011000000000000000000,
31'b0000001000000100001000000000000,
31'b0000001000000010001000000000000,
31'b0000001000000000001000000000000,
31'b0011000000100000000000000000000,
31'b0011000000100010000000000000000,
31'b0100000000000000001010010000000,
31'b0101001000000000000000000000101,
31'b0011000000101000000000000000000,
31'b0011000000101010000000000000000,
31'b0101010000010000010000000000000,
31'b0010000000000000010000010000100,
31'b0011000000110000000000000000000,
31'b0000000000000000010010000000001,
31'b0101010000001000010000000000000,
31'b0000001000101000001000000000000,
31'b0110000000000000001000000000101,
31'b0000001000100100001000000000000,
31'b0101010000000000010000000000000,
31'b0000001000100000001000000000000,
31'b0011000001000000000000000000000,
31'b0011000001000010000000000000000,
31'b0000000000000000101000000100000,
31'b0010000000001000000000000011000,
31'b0011000001001000000000000000000,
31'b0010000000000100000000000011000,
31'b0010000000000010000000000011000,
31'b0010000000000000000000000011000,
31'b0011000001010000000000000000000,
31'b0000000010000000000000000101000,
31'b0010001010000000000000100000000,
31'b0000001001001000001000000000000,
31'b0011000001011000000000000000000,
31'b0000001001000100001000000000000,
31'b0001000000000000100000100001000,
31'b0000001001000000001000000000000,
31'b0011000001100000000000000000000,
31'b0011000001100010000000000000000,
31'b0010000000000001000100010000000,
31'b1000010000000000100100000010000,
31'b0011000001101000000000000000000,
31'b1100100000000000000000100010000,
31'b1000000000000010001000011000000,
31'b1000000000000000001000011000000,
31'b1010000010000001000000000000001,
31'b0000000010100000000000000101000,
31'b0010001010100000000000100000000,
31'b0000101010000000000001000000001,
31'b1100000000000000010000001000001,
31'b0000001001100100001000000000000,
31'b0101010001000000010000000000000,
31'b0000001001100000001000000000000,
31'b0011000010000000000000000000000,
31'b0011000010000010000000000000000,
31'b0011000010000100000000000000000,
31'b0011000010000110000000000000000,
31'b0000001000000000100000000001000,
31'b0001000001000000001000100000000,
31'b0001000000010000000000000110000,
31'b0010000000000000100000100100000,
31'b0011000010010000000000000000000,
31'b0000000001000000000000000101000,
31'b0010001001000000000000100000000,
31'b0000001010001000001000000000000,
31'b0001000000000100000000000110000,
31'b0000001010000100001000000000000,
31'b0001000000000000000000000110000,
31'b0000001010000000001000000000000,
31'b1000000100000000000010000001000,
31'b1010000000000000010000000100010,
31'b1010000000000000000000111000000,
31'b1000010100000000000000001000010,
31'b0001010100000000000001000000000,
31'b0100000101000000000000001001000,
31'b0001010100000100000001000000000,
31'b0010000010000000010000010000100,
31'b1010000001000001000000000000001,
31'b0000000010000000010010000000001,
31'b0011010000000001000000001000000,
31'b0000101001000000000001000000001,
31'b0001010100010000000001000000000,
31'b0000101000000000000010001001000,
31'b0001000000100000000000000110000,
31'b0000100000000000010100000100000,
31'b0011000011000000000000000000000,
31'b0000000000010000000000000101000,
31'b0010001000010000000000100000000,
31'b0001001000000000100000000010000,
31'b0001000000000010001000100000000,
31'b0001000000000000001000100000000,
31'b0010001000011000000000100000000,
31'b0010000010000000000000000011000,
31'b0000000000000010000000000101000,
31'b0000000000000000000000000101000,
31'b0010001000000000000000100000000,
31'b0000000000000100000000000101000,
31'b0010000000000000101000000010000,
31'b0000000000001000000000000101000,
31'b0010001000001000000000100000000,
31'b0000001011000000001000000000000,
31'b1010000000010001000000000000001,
31'b0001000100000000000000000000011,
31'b0010001000110000000000100000000,
31'b0001001000100000100000000010000,
31'b0100011000000000010000100000000,
31'b0100000100000000000000001001000,
31'b1000000100000000000001001000001,
31'b1001000100000000000010000010000,
31'b1010000000000001000000000000001,
31'b0000000000100000000000000101000,
31'b0010001000100000000000100000000,
31'b0000101000000000000001000000001,
31'b1010000000001001000000000000001,
31'b0000000000101000000000000101000,
31'b0010001000101000000000100000000,
31'b0000101000001000000001000000001,
31'b0011000100000000000000000000000,
31'b1000000000010001000000000000010,
31'b1000100000000000001000001000000,
31'b1000100000000010001000001000000,
31'b1000001000000000000101000000000,
31'b1000001000000010000101000000000,
31'b1000100000001000001000001000000,
31'b0010100000000001000100000000000,
31'b1000000000000011000000000000010,
31'b1000000000000001000000000000010,
31'b1000100000010000001000001000000,
31'b1000000000000101000000000000010,
31'b1000001000010000000101000000000,
31'b1000000000001001000000000000010,
31'b0001000000000001000001001000000,
31'b0000001100000000001000000000000,
31'b1000000010000000000010000001000,
31'b1000000010000010000010000001000,
31'b1000100000100000001000001000000,
31'b1000010010000000000000001000010,
31'b0010000000000000000100000001100,
31'b0100100000000000000101000100000,
31'b0011000000000001010000000010000,
31'b0010100000100001000100000000000,
31'b1000000010010000000010000001000,
31'b1000000000100001000000000000010,
31'b1000100000000000000000000001110,
31'b1000000000000000101010000000000,
31'b0111000000000000000000001100000,
31'b1000001000000000000010100010000,
31'b0101010100000000010000000000000,
31'b0000001100100000001000000000000,
31'b1000000000000000010000000100001,
31'b1000000001010001000000000000010,
31'b0010100000000000010000000000100,
31'b0100100000001000001010000000000,
31'b1000001001000000000101000000000,
31'b0100100000000100001010000000000,
31'b0100100000000010001010000000000,
31'b0100100000000000001010000000000,
31'b1000000001000011000000000000010,
31'b1000000001000001000000000000010,
31'b0010100000010000010000000000100,
31'b1100000000000000001000010100000,
31'b1000010000000001000001000000001,
31'b1000011000000000000000000100100,
31'b0100010000000011000000000001000,
31'b0100010000000001000000000001000,
31'b1000000011000000000010000001000,
31'b0010000000000001010000000001000,
31'b0010100000100000010000000000100,
31'b0011000000000000000100000010100,
31'b0100110000010000000000000000100,
31'b0100000010000000000000001001000,
31'b1000001000000000001010000100000,
31'b1001000010000000000010000010000,
31'b0100110000001000000000000000100,
31'b1011000000000000000010000100000,
31'b0000101000000000001000010000000,
31'b1001000000000000000100010000010,
31'b0100110000000000000000000000100,
31'b0100110000000010000000000000100,
31'b0100000000000000101000001000000,
31'b0100010000100001000000000001000,
31'b1000000000100000000010000001000,
31'b1000000010010001000000000000010,
31'b1000100010000000001000001000000,
31'b1000100000000001000010000000100,
31'b0001010000100000000001000000000,
31'b0100001000000000011001000000000,
31'b0001010000100100000001000000000,
31'b0010100010000001000100000000000,
31'b1000000010000011000000000000010,
31'b1000000010000001000000000000010,
31'b0111000000000000010001000000000,
31'b1000010000000000001000000001100,
31'b0001010000110000000001000000000,
31'b1100001000000000000000010001000,
31'b0001000100000000000000000110000,
31'b0000001110000000001000000000000,
31'b1000000000000000000010000001000,
31'b1000000000000010000010000001000,
31'b1000000000000100000010000001000,
31'b1000010000000000000000001000010,
31'b0001010000000000000001000000000,
31'b0100000001000000000000001001000,
31'b0001010000000100000001000000000,
31'b1001000001000000000010000010000,
31'b1000000000010000000010000001000,
31'b1000000010100001000000000000010,
31'b1000000000010100000010000001000,
31'b1000010000010000000000001000010,
31'b0001010000010000000001000000000,
31'b0110000000000000000001010000100,
31'b0001010000010100000001000000000,
31'b0010101000000000000000110000000,
31'b1000000010000000010000000100001,
31'b0001000000100000000000000000011,
31'b0010100010000000010000000000100,
31'b0001001100000000100000000010000,
31'b0100010000000001101000000000000,
31'b0100000000100000000000001001000,
31'b1000100000000000010110000000000,
31'b1010100000000000000000101000000,
31'b0010000000000000010010000000010,
31'b0000000100000000000000000101000,
31'b0010001100000000000000100000000,
31'b0000011000000000000000010000010,
31'b0100100000000000100010000001000,
31'b0100000000000000001000000000110,
31'b1010000000000000010000000010001,
31'b0100010010000001000000000001000,
31'b1000000001000000000010000001000,
31'b0001000000000000000000000000011,
31'b1000000001000100000010000001000,
31'b0001000000000100000000000000011,
31'b0100000000000010000000001001000,
31'b0100000000000000000000001001000,
31'b1000000000000000000001001000001,
31'b1001000000000000000010000010000,
31'b1010000100000001000000000000001,
31'b0001000000010000000000000000011,
31'b0010001100100000000000100000000,
31'b0001100000000000000000010110000,
31'b0100110010000000000000000000100,
31'b0100000000010000000000001001000,
31'b1010000000000000100010100000000,
31'b1001000000010000000010000010000,
31'b0011001000000000000000000000000,
31'b0011001000000010000000000000000,
31'b0011001000000100000000000000000,
31'b0000000000011000001000000000000,
31'b0000000010000000100000000001000,
31'b0000000000010100001000000000000,
31'b0000000000010010001000000000000,
31'b0000000000010000001000000000000,
31'b0011001000010000000000000000000,
31'b0000000000001100001000000000000,
31'b0000000000001010001000000000000,
31'b0000000000001000001000000000000,
31'b0000000000000110001000000000000,
31'b0000000000000100001000000000000,
31'b0000000000000010001000000000000,
31'b0000000000000000001000000000000,
31'b0011001000100000000000000000000,
31'b0110010000000000011000000000000,
31'b0101000000000010000000000000101,
31'b0101000000000000000000000000101,
31'b0000010000000000000010000000100,
31'b0000010000000010000010000000100,
31'b0000010000000100000010000000100,
31'b0000000000110000001000000000000,
31'b0011001000110000000000000000000,
31'b0000001000000000010010000000001,
31'b0010010000000000000000010000001,
31'b0000000000101000001000000000000,
31'b0000010000010000000010000000100,
31'b0000000000100100001000000000000,
31'b0000000000100010001000000000000,
31'b0000000000100000001000000000000,
31'b0011001001000000000000000000000,
31'b0011001001000010000000000000000,
31'b0010000010010000000000100000000,
31'b0001000010000000100000000010000,
31'b0000000000000000000000100110000,
31'b0000000001010100001000000000000,
31'b0000000001010010001000000000000,
31'b0000000001010000001000000000000,
31'b0010000010000100000000100000000,
31'b0000001010000000000000000101000,
31'b0010000010000000000000100000000,
31'b0000000001001000001000000000000,
31'b0000000001000110001000000000000,
31'b0000000001000100001000000000000,
31'b0000000001000010001000000000000,
31'b0000000001000000001000000000000,
31'b0011001001100000000000000000000,
31'b1100010000000000000000001000100,
31'b0010001000000001000100010000000,
31'b1100100000000000101000000000000,
31'b0000010001000000000010000000100,
31'b1000010000000000001100100000000,
31'b1000000100000000001010000100000,
31'b1000000000000000000001000010100,
31'b1100100010000000000000000001000,
31'b0000100010000100000001000000001,
31'b0010000010100000000000100000000,
31'b0000100010000000000001000000001,
31'b0000010100000100000001100000000,
31'b0000000001100100001000000000000,
31'b0000010100000000000001100000000,
31'b0000000001100000001000000000000,
31'b0000000000001000100000000001000,
31'b0010000000000000001000000110000,
31'b0010000001010000000000100000000,
31'b0001000001000000100000000010000,
31'b0000000000000000100000000001000,
31'b0000000000000010100000000001000,
31'b0000000000000100100000000001000,
31'b0000000010010000001000000000000,
31'b0010000001000100000000100000000,
31'b0000001001000000000000000101000,
31'b0010000001000000000000100000000,
31'b0000000010001000001000000000000,
31'b0000000000010000100000000001000,
31'b0000000010000100001000000000000,
31'b0000000010000010001000000000000,
31'b0000000010000000001000000000000,
31'b1010010000000000000100000000000,
31'b1010010000000010000100000000000,
31'b1010010000000100000100000000000,
31'b0101000010000000000000000000101,
31'b0000000000100000100000000001000,
31'b0000010000000001001000001000000,
31'b0000110000010000000000000000010,
31'b0000100000000001100000000000100,
31'b1100100001000000000000000001000,
31'b0000100001000100000001000000001,
31'b0010000001100000000000100000000,
31'b0000100001000000000001000000001,
31'b0000110000000100000000000000010,
31'b0000100000000000000010001001000,
31'b0000110000000000000000000000010,
31'b0000000010100000001000000000000,
31'b0010000000010100000000100000000,
31'b0001000000000100100000000010000,
31'b0010000000010000000000100000000,
31'b0001000000000000100000000010000,
31'b0000000001000000100000000001000,
31'b0001001000000000001000100000000,
31'b0010000000011000000000100000000,
31'b0001000000001000100000000010000,
31'b0010000000000100000000100000000,
31'b0000001000000000000000000101000,
31'b0010000000000000000000100000000,
31'b0010000000000010000000100000000,
31'b0010000000001100000000100000000,
31'b0000001000001000000000000101000,
31'b0010000000001000000000100000000,
31'b0000000011000000001000000000000,
31'b1100100000010000000000000001000,
31'b0001001100000000000000000000011,
31'b0010000000110000000000100000000,
31'b0001000000100000100000000010000,
31'b0100010000000000010000100000000,
31'b0100010000000010010000100000000,
31'b0110000000000000000100000001010,
31'b1001000000000001001000000000001,
31'b1100100000000000000000000001000,
31'b0000100000000100000001000000001,
31'b0010000000100000000000100000000,
31'b0000100000000000000001000000001,
31'b1100100000001000000000000001000,
31'b0000100001000000000010001001000,
31'b0010000000101000000000100000000,
31'b0000100000001000000001000000001,
31'b1000000000001000000101000000000,
31'b1000001000010001000000000000010,
31'b1000101000000000001000001000000,
31'b0001000000000000000100001000010,
31'b1000000000000000000101000000000,
31'b1000000000000010000101000000000,
31'b1000000000000100000101000000000,
31'b0000000100010000001000000000000,
31'b1000001000000011000000000000010,
31'b1000001000000001000000000000010,
31'b0010100000000000000001000000010,
31'b0000000100001000001000000000000,
31'b1000000000010000000101000000000,
31'b0000000100000100001000000000000,
31'b0000000100000010001000000000000,
31'b0000000100000000001000000000000,
31'b1000001010000000000010000001000,
31'b0100100001000000010000000000001,
31'b0100000000000010001000001100000,
31'b0100000000000000001000001100000,
31'b1000000000100000000101000000000,
31'b1000000000100010000101000000000,
31'b1000000001000000001010000100000,
31'b0000000100110000001000000000000,
31'b0100100000000001000000000100010,
31'b0000000000000100000000100000011,
31'b0000100001000000001000010000000,
31'b0000000000000000000000100000011,
31'b1000000000110000000101000000000,
31'b1000000000000000000010100010000,
31'b0000010001000000000001100000000,
31'b0000000100100000001000000000000,
31'b1000001000000000010000000100001,
31'b1000010000000000000100000000011,
31'b0010101000000000010000000000100,
31'b0001000110000000100000000010000,
31'b1000000001000000000101000000000,
31'b1000010000010000000000000100100,
31'b1000000001000100000101000000000,
31'b0000010000000000000110000010000,
31'b0111100000000000000010000000000,
31'b1000010000001000000000000100100,
31'b0010000110000000000000100000000,
31'b0000010010000000000000010000010,
31'b1000010000000010000000000100100,
31'b1000010000000000000000000100100,
31'b0000010000100000000001100000000,
31'b0000000101000000001000000000000,
31'b0100100000000010010000000000001,
31'b0100100000000000010000000000001,
31'b0000100000010000001000010000000,
31'b0100100000000100010000000000001,
31'b1000000001100000000101000000000,
31'b0100100000001000010000000000001,
31'b1000000000000000001010000100000,
31'b1000000100000000000001000010100,
31'b0100000000000000000000101010000,
31'b0100100000010000010000000000001,
31'b0000100000000000001000010000000,
31'b0000100000000010001000010000000,
31'b0000010000000100000001100000000,
31'b1000010000100000000000000100100,
31'b0000010000000000000001100000000,
31'b0000010000000010000001100000000,
31'b0010000000000000000011000000100,
31'b0100100000000000000010000101000,
31'b0010000101010000000000100000000,
31'b0001000101000000100000000010000,
31'b0000000100000000100000000001000,
31'b0100000000000000011001000000000,
31'b0000000100000100100000000001000,
31'b0000000110010000001000000000000,
31'b0010000101000100000000100000000,
31'b1100000000001000000000010001000,
31'b0010000101000000000000100000000,
31'b0000010001000000000000010000010,
31'b0000000100010000100000000001000,
31'b1100000000000000000000010001000,
31'b0000000000000000000001010000001,
31'b0000000110000000001000000000000,
31'b1000001000000000000010000001000,
31'b1000001000000010000010000001000,
31'b1000001000000100000010000001000,
31'b1010000000000000000010100100000,
31'b0001011000000000000001000000000,
31'b0100001001000000000000001001000,
31'b0001100000000000100000010010000,
31'b0010100000010000000000110000000,
31'b1100000000000001000100000010000,
31'b0010010000000100001001000000000,
31'b0010010000000010001001000000000,
31'b0010010000000000001001000000000,
31'b0001011000010000000001000000000,
31'b1100000000100000000000010001000,
31'b0000110100000000000000000000010,
31'b0010100000000000000000110000000,
31'b0010000100010100000000100000000,
31'b0001001000100000000000000000011,
31'b0010000100010000000000100000000,
31'b0001000100000000100000000010000,
31'b0000000101000000100000000001000,
31'b0100001000100000000000001001000,
31'b0010000100011000000000100000000,
31'b0001000100001000100000000010000,
31'b0010000100000100000000100000000,
31'b0000010000000100000000010000010,
31'b0010000100000000000000100000000,
31'b0000010000000000000000010000010,
31'b0010000100001100000000100000000,
31'b1100000001000000000000010001000,
31'b0010000100001000000000100000000,
31'b0000010000001000000000010000010,
31'b1000100000000000001100000000001,
31'b0001001000000000000000000000011,
31'b0010000100110000000000100000000,
31'b0001001000000100000000000000011,
31'b0100010100000000010000100000000,
31'b0100001000000000000000001001000,
31'b1000001000000000000001001000001,
31'b1001001000000000000010000010000,
31'b1100100100000000000000000001000,
31'b0001010000000000100001000100000,
31'b0010000100100000000000100000000,
31'b0000100100000000000001000000001,
31'b0010000000000100001000000000011,
31'b1100000000000000010000000010100,
31'b0010000000000000001000000000011,
31'b0010100001000000000000110000000,
31'b0011010000000000000000000000000,
31'b0100000000010000000000010000100,
31'b0011010000000100000000000000000,
31'b0110000000001000000010000000001,
31'b0011010000001000000000000000000,
31'b0110000000000100000010000000001,
31'b0110000000000010000010000000001,
31'b0110000000000000000010000000001,
31'b0100000000000010000000010000100,
31'b0100000000000000000000010000100,
31'b0101000000101000010000000000000,
31'b0100000000000100000000010000100,
31'b0101000000100100010000000000000,
31'b0100000000001000000000010000100,
31'b0101000000100000010000000000000,
31'b0000011000000000001000000000000,
31'b0011010000100000000000000000000,
31'b0110001000000000011000000000000,
31'b0101000000011000010000000000000,
31'b1000000110000000000000001000010,
31'b0000001000000000000010000000100,
31'b0001000000000000001000010000001,
31'b0101000000010000010000000000000,
31'b0110000000100000000010000000001,
31'b0101000000001100010000000000000,
31'b0100000000100000000000010000100,
31'b0101000000001000010000000000000,
31'b0101000000001010010000000000000,
31'b0101000000000100010000000000000,
31'b0101000000000110010000000000000,
31'b0101000000000000010000000000000,
31'b0101000000000010010000000000000,
31'b0011010001000000000000000000000,
31'b0110000000000000000001001001000,
31'b1010000000000000000000001000001,
31'b1010000000000010000000001000001,
31'b0011010001001000000000000000000,
31'b0011000000000000000001000000011,
31'b1010000000001000000000001000001,
31'b0010010000000000000000000011000,
31'b0101100000000000000100000001000,
31'b0100000001000000000000010000100,
31'b1010000000010000000000001000001,
31'b0100000100001001000000000001000,
31'b1000000100000001000001000000001,
31'b1000001100000000000000000100100,
31'b0101000001100000010000000000000,
31'b0100000100000001000000000001000,
31'b0011010001100000000000000000000,
31'b1100001000000000000000001000100,
31'b1010000000100000000000001000001,
31'b1000000000000000100100000010000,
31'b0001100000000000000000100000010,
31'b1000100000000000100000010000100,
31'b0101000001010000010000000000000,
31'b1000010000000000001000011000000,
31'b0100100100001000000000000000100,
31'b0100000000000000010000000011000,
31'b1011000000000000000100100000000,
31'b1001000000000000010010001000000,
31'b0100100100000000000000000000100,
31'b0100100100000010000000000000100,
31'b0101000001000000010000000000000,
31'b0101000001000010010000000000000,
31'b0011010010000000000000000000000,
31'b0110100000000000000100000100000,
31'b0011010010000100000000000000000,
31'b1100000000000000000100000000101,
31'b0001000100100000000001000000000,
31'b0001010001000000001000100000000,
31'b0001010000010000000000000110000,
31'b1100000000010000000000000100010,
31'b0101000000000000000001001100000,
31'b0100000010000000000000010000100,
31'b0011000000100001000000001000000,
31'b1100000000001000000000000100010,
31'b0001010000000100000000000110000,
31'b1100000000000100000000000100010,
31'b0001010000000000000000000110000,
31'b1100000000000000000000000100010,
31'b1010001000000000000100000000000,
31'b1010001000000010000100000000000,
31'b1010001000000100000100000000000,
31'b1000000100000000000000001000010,
31'b0001000100000000000001000000000,
31'b0001000100000010000001000000000,
31'b0001000100000100000001000000000,
31'b1001000000010000001100000000000,
31'b1010001000010000000100000000000,
31'b0100000010100000000000010000100,
31'b0011000000000001000000001000000,
31'b1001000000001000001100000000000,
31'b0001000100010000000001000000000,
31'b1010000000000001000001000000010,
31'b0000101000000000000000000000010,
31'b1001000000000000001100000000000,
31'b0011010011000000000000000000000,
31'b0001100000000000000001010000000,
31'b1100001000000000100000000000010,
31'b0001100000000100000001010000000,
31'b0100001000100000010000100000000,
31'b0001010000000000001000100000000,
31'b1100000000000001010000000000001,
31'b0010010010000000000000000011000,
31'b0010000000000000000100011000000,
31'b0000010000000000000000000101000,
31'b0010011000000000000000100000000,
31'b0000010000000100000000000101000,
31'b1000000000000011001000010000000,
31'b1000000000000001001000010000000,
31'b0010100000000000000000001010100,
31'b1100000001000000000000000100010,
31'b1100000100000000000000000010001,
31'b0001100000100000000001010000000,
31'b0100000100001000000010000000010,
31'b0000100000000000100000000100010,
31'b0100001000000000010000100000000,
31'b0100010100000000000000001001000,
31'b0100000100000000000010000000010,
31'b0110000000000000010000000101000,
31'b1010010000000001000000000000001,
31'b0000010000100000000000000101000,
31'b0011000001000001000000001000000,
31'b0000111000000000000001000000001,
31'b0100100110000000000000000000100,
31'b1010000000000000100100000100000,
31'b0001000000000000000010100000100,
31'b1001000001000000001100000000000,
31'b1000000000000000100000000000100,
31'b1000000000000010100000000000100,
31'b1000000000000100100000000000100,
31'b1000000010100000000000001000010,
31'b1000000000001000100000000000100,
31'b1000000000001010100000000000100,
31'b1000000000001100100000000000100,
31'b0110000100000000000010000000001,
31'b1000000000010000100000000000100,
31'b1000010000000001000000000000010,
31'b1000000000010100100000000000100,
31'b1000010000000101000000000000010,
31'b1000000001000001000001000000001,
31'b1000010000001001000000000000010,
31'b0101000100100000010000000000000,
31'b0100000001000001000000000001000,
31'b1000000000100000100000000000100,
31'b1000000010000100000000001000010,
31'b1000000010000010000000001000010,
31'b1000000010000000000000001000010,
31'b0001000010000000000001000000000,
31'b0001000010000010000001000000000,
31'b0001000010000100000001000000000,
31'b1001000000000000110000010000000,
31'b1000100010000001001000000000000,
31'b1000100000000000000010001000100,
31'b0101000100001000010000000000000,
31'b1000010000000000101010000000000,
31'b0100100001000000000000000000100,
31'b0101000000000000000100010001000,
31'b0101000100000000010000000000000,
31'b0101000100000010010000000000000,
31'b1000000001000000100000000000100,
31'b1000001000000000000100000000011,
31'b1010000100000000000000001000001,
31'b0100000000011001000000000001000,
31'b1000000001001000100000000000100,
31'b1000001000010000000000000100100,
31'b0100000010100000000010000000010,
31'b0100000000010001000000000001000,
31'b1000000001010000100000000000100,
31'b1000010001000001000000000000010,
31'b0100000000100000000100010010000,
31'b0100000000001001000000000001000,
31'b1000000000000001000001000000001,
31'b1000001000000000000000000100100,
31'b0100000000000011000000000001000,
31'b0100000000000001000000000001000,
31'b1100000010000000000000000010001,
31'b0011000000000000001001100000000,
31'b0100000010001000000010000000010,
31'b0000000010000000000001000011000,
31'b0100100000010000000000000000100,
31'b0100100000010010000000000000100,
31'b0100000010000000000010000000010,
31'b0100000010000010000010000000010,
31'b0100100000001000000000000000100,
31'b0100100000001010000000000000100,
31'b0100000000000000000100010010000,
31'b0100000000101001000000000001000,
31'b0100100000000000000000000000100,
31'b0100100000000010000000000000100,
31'b0000001000000000000001100000000,
31'b0100000000100001000000000001000,
31'b1000000010000000100000000000100,
31'b1000000010000010100000000000100,
31'b1000000010000100100000000000100,
31'b1000000000100000000000001000010,
31'b0001000000100000000001000000000,
31'b0001000000100010000001000000000,
31'b0001000000100100000001000000000,
31'b1001000000000000000000100100100,
31'b1000100000100001001000000000000,
31'b1000010010000001000000000000010,
31'b1000100000000000100010000000010,
31'b1000000000000000001000000001100,
31'b0001000000110000000001000000000,
31'b0010100000100000000100001000000,
31'b0001010100000000000000000110000,
31'b1100000100000000000000000100010,
31'b0001000000001000000001000000000,
31'b1000000000000100000000001000010,
31'b1000000000000010000000001000010,
31'b1000000000000000000000001000010,
31'b0001000000000000000001000000000,
31'b0001000000000010000001000000000,
31'b0001000000000100000001000000000,
31'b1000000000001000000000001000010,
31'b1000100000000001001000000000000,
31'b1000100000000011001000000000000,
31'b1000100000000101001000000000000,
31'b1000000000010000000000001000010,
31'b0001000000010000000001000000000,
31'b0010100000000000000100001000000,
31'b0001000000010100000001000000000,
31'b1001000100000000001100000000000,
31'b1100000000100000000000000010001,
31'b0001100100000000000001010000000,
31'b0100001000000001000000100010000,
31'b0000001000010000000000010000010,
31'b0100000000000001101000000000000,
31'b0100010000100000000000001001000,
31'b0100000000100000000010000000010,
31'b0100000010010001000000000001000,
31'b0010010000000000010010000000010,
31'b0000010100000000000000000101000,
31'b0000001000000010000000010000010,
31'b0000001000000000000000010000010,
31'b1001000000000000001000000010100,
31'b1000001010000000000000000100100,
31'b0100000010000011000000000001000,
31'b0100000010000001000000000001000,
31'b1100000000000000000000000010001,
31'b0001010000000000000000000000011,
31'b0100000000001000000010000000010,
31'b0000000000000000000001000011000,
31'b0001000001000000000001000000000,
31'b0100010000000000000000001001000,
31'b0100000000000000000010000000010,
31'b0100000000000010000010000000010,
31'b1100000000010000000000000010001,
31'b0001010000010000000000000000011,
31'b0100000010000000000100010010000,
31'b0000001000100000000000010000010,
31'b0100100010000000000000000000100,
31'b0100100010000010000000000000100,
31'b0100000000010000000010000000010,
31'b0100000010100001000000000001000,
31'b0011011000000000000000000000000,
31'b0110000000100000011000000000000,
31'b0011011000000100000000000000000,
31'b0001000000000000010010010000000,
31'b0000000000100000000010000000100,
31'b0000010000010100001000000000000,
31'b0000010000010010001000000000000,
31'b0000010000010000001000000000000,
31'b0101000000000000001010000000001,
31'b0100001000000000000000010000100,
31'b0010000000100000000000010000001,
31'b0000010000001000001000000000000,
31'b0000010000000110001000000000000,
31'b0000010000000100001000000000000,
31'b0000010000000010001000000000000,
31'b0000010000000000001000000000000,
31'b0000000000001000000010000000100,
31'b0110000000000000011000000000000,
31'b0010000000010000000000010000001,
31'b0110000000000100011000000000000,
31'b0000000000000000000010000000100,
31'b0000000000000010000010000000100,
31'b0000000000000100000010000000100,
31'b0000010000110000001000000000000,
31'b0010000000000100000000010000001,
31'b0110000000010000011000000000000,
31'b0010000000000000000000010000001,
31'b0010000000000010000000010000001,
31'b0000000000010000000010000000100,
31'b0000010000100100001000000000000,
31'b0000100010000000000000000000010,
31'b0000010000100000001000000000000,
31'b0011011001000000000000000000000,
31'b1100000000100000000000001000100,
31'b1100000010000000100000000000010,
31'b0001010010000000100000000010000,
31'b0000010000000000000000100110000,
31'b1000000100010000000000000100100,
31'b0000010001010010001000000000000,
31'b0000010001010000001000000000000,
31'b0011000000000001000100000000001,
31'b1100000000000000001000000001010,
31'b0010010010000000000000100000000,
31'b0000010001001000001000000000000,
31'b1000000100000010000000000100100,
31'b1000000100000000000000000100100,
31'b0000010001000010001000000000000,
31'b0000010001000000001000000000000,
31'b0010000000000001000000101000000,
31'b1100000000000000000000001000100,
31'b0010000001010000000000010000001,
31'b1100000000000100000000001000100,
31'b0000000001000000000010000000100,
31'b1000000000000000001100100000000,
31'b0000000100010000000001100000000,
31'b1000010000000000000001000010100,
31'b0010000001000100000000010000001,
31'b1100000000010000000000001000100,
31'b0010000001000000000000010000001,
31'b0010100000000000001000100000010,
31'b0000000100000100000001100000000,
31'b1000000100100000000000000100100,
31'b0000000100000000000001100000000,
31'b0000010001100000001000000000000,
31'b1010000000100000000100000000000,
31'b1010000000100010000100000000000,
31'b1100000001000000100000000000010,
31'b0001010001000000100000000010000,
31'b0000010000000000100000000001000,
31'b0000010000000010100000000001000,
31'b0000100000110000000000000000010,
31'b0000010010010000001000000000000,
31'b1010000000110000000100000000000,
31'b0100001010000000000000010000100,
31'b0010010001000000000000100000000,
31'b0000010010001000001000000000000,
31'b0000100000100100000000000000010,
31'b0000010010000100001000000000000,
31'b0000100000100000000000000000010,
31'b0000010010000000001000000000000,
31'b1010000000000000000100000000000,
31'b1010000000000010000100000000000,
31'b1010000000000100000100000000000,
31'b1010000000000110000100000000000,
31'b0000000010000000000010000000100,
31'b0000000000000001001000001000000,
31'b0000100000010000000000000000010,
31'b0000100000010010000000000000010,
31'b1010000000010000000100000000000,
31'b1010000000010010000100000000000,
31'b0000100000001000000000000000010,
31'b0010000100000000001001000000000,
31'b0000100000000100000000000000010,
31'b0000100000000110000000000000010,
31'b0000100000000000000000000000010,
31'b0000100000000010000000000000010,
31'b1100000000000100100000000000010,
31'b0001101000000000000001010000000,
31'b1100000000000000100000000000010,
31'b0001010000000000100000000010000,
31'b0100000000100000010000100000000,
31'b0101000000000000100001001000000,
31'b1100000000001000100000000000010,
31'b0001010000001000100000000010000,
31'b0010010000000100000000100000000,
31'b0000011000000000000000000101000,
31'b0010010000000000000000100000000,
31'b0000000100000000000000010000010,
31'b0110100000000000100100000000000,
31'b1000001000000001001000010000000,
31'b0010010000001000000000100000000,
31'b0000010011000000001000000000000,
31'b1010000001000000000100000000000,
31'b1100000010000000000000001000100,
31'b1100000000100000100000000000010,
31'b0001010000100000100000000010000,
31'b0100000000000000010000100000000,
31'b0100000000000010010000100000000,
31'b0100000000000100010000100000000,
31'b0100000000000110010000100000000,
31'b1100110000000000000000000001000,
31'b0001100000000000000000000011010,
31'b0010010000100000000000100000000,
31'b0000110000000000000001000000001,
31'b0100000000010000010000100000000,
31'b0100100000000000000000001010001,
31'b0000100001000000000000000000010,
31'b0000100001000010000000000000010,
31'b1000001000000000100000000000100,
31'b1000001000000010100000000000100,
31'b1100000000000000000100001010000,
31'b0001010000000000000100001000010,
31'b1000010000000000000101000000000,
31'b1000010000000010000101000000000,
31'b1000010000000100000101000000000,
31'b0000010100010000001000000000000,
31'b1000001000010000100000000000100,
31'b1000011000000001000000000000010,
31'b0010110000000000000001000000010,
31'b0000010100001000001000000000000,
31'b1000010000010000000101000000000,
31'b1000000001000000000000000100100,
31'b0000010100000010001000000000000,
31'b0000010100000000001000000000000,
31'b0010000000000000100001000001000,
31'b0110000100000000011000000000000,
31'b0010000100010000000000010000001,
31'b1110000000000000100000000000001,
31'b0000000100000000000010000000100,
31'b0000000100000010000010000000100,
31'b0000000100000100000010000000100,
31'b0000010100110000001000000000000,
31'b0010000100000100000000010000001,
31'b0010000010000100001001000000000,
31'b0010000100000000000000010000001,
31'b0010000010000000001001000000000,
31'b0000000100010000000010000000100,
31'b1000010000000000000010100010000,
31'b0000000001000000000001100000000,
31'b0000010100100000001000000000000,
31'b1000001001000000100000000000100,
31'b1000000000000000000100000000011,
31'b0100000010000001000000100010000,
31'b0000000010010000000000010000010,
31'b1000010001000000000101000000000,
31'b1000000000010000000000000100100,
31'b0000000000110000000001100000000,
31'b0000000000000000000110000010000,
31'b1000000000001010000000000100100,
31'b1000000000001000000000000100100,
31'b0000000010000010000000010000010,
31'b0000000010000000000000010000010,
31'b1000000000000010000000000100100,
31'b1000000000000000000000000100100,
31'b0000000000100000000001100000000,
31'b0010100000000000000000000000001,
31'b0010000100000001000000101000000,
31'b1100000100000000000000001000100,
31'b0000000000011000000001100000000,
31'b0000001010000000000001000011000,
31'b0000000101000000000010000000100,
31'b1000000100000000001100100000000,
31'b0000000000010000000001100000000,
31'b0000000000100000000110000010000,
31'b0000000000001100000001100000000,
31'b1001000000000000000000101000010,
31'b0000000000001000000001100000000,
31'b0000000010100000000000010000010,
31'b0000000000000100000001100000000,
31'b1000000000100000000000000100100,
31'b0000000000000000000001100000000,
31'b0000000000000010000001100000000,
31'b1010000100100000000100000000000,
31'b0100100000000000010000110000000,
31'b0100100000000000000000001100010,
31'b0000000001010000000000010000010,
31'b0001001000100000000001000000000,
31'b0101000000000001000000100001000,
31'b0001100000000000000000000101001,
31'b0000010110010000001000000000000,
31'b0100000000000011001000000100000,
31'b0100000000000001001000000100000,
31'b0000100000000000001000100000001,
31'b0000000001000000000000010000010,
31'b0001001000110000000001000000000,
31'b1100010000000000000000010001000,
31'b0000100100100000000000000000010,
31'b0000010110000000001000000000000,
31'b1010000100000000000100000000000,
31'b1010000100000010000100000000000,
31'b1010000100000100000100000000000,
31'b1000001000000000000000001000010,
31'b0001001000000000000001000000000,
31'b0001001000000010000001000000000,
31'b0001001000000100000001000000000,
31'b1011100000000001000000000000000,
31'b1010000100010000000100000000000,
31'b0010000000000100001001000000000,
31'b0010000000000010001001000000000,
31'b0010000000000000001001000000000,
31'b0001001000010000000001000000000,
31'b0010101000000000000100001000000,
31'b0000100100000000000000000000010,
31'b0010000000001000001001000000000,
31'b0100000000000101000000100010000,
31'b0000100000000000000000000110001,
31'b0100000000000001000000100010000,
31'b0000000000010000000000010000010,
31'b0100001000000001101000000000000,
31'b1010100000000000000100010000000,
31'b0100001000100000000010000000010,
31'b0000000010000000000110000010000,
31'b0000000000000110000000010000010,
31'b0000000000000100000000010000010,
31'b0000000000000010000000010000010,
31'b0000000000000000000000010000010,
31'b1001000000000000000001011000000,
31'b1000000010000000000000000100100,
31'b0000000010100000000001100000000,
31'b0000000000001000000000010000010,
31'b1100001000000000000000000010001,
31'b0001011000000000000000000000011,
31'b0100001000001000000010000000010,
31'b0000001000000000000001000011000,
31'b0100000100000000010000100000000,
31'b0100011000000000000000001001000,
31'b0100001000000000000010000000010,
31'b0100001000000010000010000000010,
31'b0001000000001000010000000000110,
31'b0001000000000000100001000100000,
31'b0000000010001000000001100000000,
31'b0000000000100000000000010000010,
31'b0001000000000000010000000000110,
31'b1000000010100000000000000100100,
31'b0000000010000000000001100000000,
31'b0000000010000010000001100000000,
31'b0011100000000000000000000000000,
31'b0011100000000010000000000000000,
31'b1000000100000000001000001000000,
31'b1001001000000001000001000000000,
31'b0011100000001000000000000000000,
31'b0011100000001010000000000000000,
31'b1001000000010000000100000000010,
31'b0010000100000001000100000000000,
31'b0011100000010000000000000000000,
31'b0000000000000000000101001000000,
31'b1001000000001000000100000000010,
31'b0000101000001000001000000000000,
31'b1010000000000001001001000000000,
31'b0000101000000100001000000000000,
31'b1001000000000000000100000000010,
31'b0000101000000000001000000000000,
31'b0011100000100000000000000000000,
31'b0010000000000000010100000010000,
31'b1101000000000000000000100001000,
31'b0011000000000001000000000001100,
31'b0011100000101000000000000000000,
31'b1100000001000000000000100010000,
31'b1100000000010000001000000100000,
31'b0010100000000000010000010000100,
31'b0011100000110000000000000000000,
31'b0000100000000000010010000000001,
31'b1100000000001000001000000100000,
31'b0000101000101000001000000000000,
31'b1100000000000100001000000100000,
31'b0000101000100100001000000000000,
31'b1100000000000000001000000100000,
31'b0000101000100000001000000000000,
31'b0011100001000000000000000000000,
31'b0011100001000010000000000000000,
31'b0010000100000000010000000000100,
31'b0100000100001000001010000000000,
31'b0011100001001000000000000000000,
31'b1100000000100000000000100010000,
31'b0100000100000010001010000000000,
31'b0100000100000000001010000000000,
31'b0110000010000000000001000000100,
31'b0000100010000000000000000101000,
31'b0010101010000000000000100000000,
31'b0000101001001000001000000000000,
31'b1100000000000000000111000000000,
31'b0000101001000100001000000000000,
31'b1001000001000000000100000000010,
31'b0000101001000000001000000000000,
31'b0011100001100000000000000000000,
31'b1100000000001000000000100010000,
31'b0010100000000001000100010000000,
31'b1100001000000000101000000000000,
31'b0010000000000001000000000010100,
31'b1100000000000000000000100010000,
31'b0011000000000000010100000001000,
31'b1100000000000100000000100010000,
31'b1100001010000000000000000001000,
31'b0000100010100000000000000101000,
31'b0000001100000000001000010000000,
31'b0000001010000000000001000000001,
31'b1000000000000001000000010000010,
31'b1100000000010000000000100010000,
31'b1100000001000000001000000100000,
31'b0000101001100000001000000000000,
31'b0100000000000000000000011001000,
31'b0110010000000000000100000100000,
31'b1001000000000000000010010010000,
31'b1000000100000001000010000000100,
31'b0001000000000000000000010000011,
31'b1000000001000000000010010001000,
31'b0001100000010000000000000110000,
31'b0010100000000000100000100100000,
31'b0110000001000000000001000000100,
31'b0000100001000000000000000101000,
31'b0011000000000000000010000000110,
31'b0000101010001000001000000000000,
31'b0001100000000100000000000110000,
31'b0000101010000100001000000000000,
31'b0001100000000000000000000110000,
31'b0000101010000000001000000000000,
31'b1110000000000000001000000010000,
31'b0011010000000000001000000000010,
31'b0000011000011000000000000000010,
31'b0000010000000001000101000000000,
31'b0001110100000000000001000000000,
31'b1100000000000000100000000101000,
31'b0000011000010000000000000000010,
31'b0000001000000001100000000000100,
31'b1100001001000000000000000001000,
31'b0000100010000000010010000000001,
31'b0000011000001000000000000000010,
31'b0000001001000000000001000000001,
31'b0000011000000100000000000000010,
31'b0000001000000000000010001001000,
31'b0000011000000000000000000000010,
31'b0000000000000000010100000100000,
31'b0110000000010000000001000000100,
31'b0001010000000000000001010000000,
31'b0010101000010000000000100000000,
31'b0001101000000000100000000010000,
31'b1000001000000000000100100000010,
31'b1000000000000000000010010001000,
31'b1000010000000000000000011000010,
31'b1010000100000000000000101000000,
31'b0110000000000000000001000000100,
31'b0000100000000000000000000101000,
31'b0010101000000000000000100000000,
31'b0000100000000100000000000101000,
31'b0110000000001000000001000000100,
31'b0000100000001000000000000101000,
31'b0010101000001000000000100000000,
31'b0000101011000000001000000000000,
31'b1100001000010000000000000001000,
31'b0001100100000000000000000000011,
31'b0000001000000000110100000000000,
31'b0000010000000000100000000100010,
31'b0011000000000000001001000000001,
31'b1100000010000000000000100010000,
31'b0000010000000000010001000000100,
31'b0000010000001000100000000100010,
31'b1100001000000000000000000001000,
31'b0000100000100000000000000101000,
31'b0000000000000001000000000100100,
31'b0000001000000000000001000000001,
31'b1100001000001000000000000001000,
31'b0000100000101000000000000101000,
31'b0000011001000000000000000000010,
31'b0000001000001000000001000000001,
31'b1000000000000100001000001000000,
31'b1000100000010001000000000000010,
31'b1000000000000000001000001000000,
31'b1000000000000010001000001000000,
31'b1000101000000000000101000000000,
31'b0010000000000101000100000000000,
31'b1000000000001000001000001000000,
31'b0010000000000001000100000000000,
31'b1000100000000011000000000000010,
31'b1000100000000001000000000000010,
31'b1000000000010000001000001000000,
31'b1000100000000101000000000000010,
31'b0100010001100000000000000000100,
31'b1011001000000000000000001000000,
31'b1001000100000000000100000000010,
31'b0010000000010001000100000000000,
31'b1000100010000000000010000001000,
31'b0100001001000000010000000000001,
31'b1000000000100000001000001000000,
31'b1000010000000001100000000001000,
31'b0100010001010000000000000000100,
31'b0100000000000000000101000100000,
31'b1000000000101000001000001000000,
31'b0010000000100001000100000000000,
31'b1000010010000001001000000000000,
31'b1000100000100001000000000000010,
31'b1000000000000000000000000001110,
31'b1000100000000000101010000000000,
31'b0100010001000000000000000000100,
31'b0100010001000010000000000000100,
31'b1100000100000000001000000100000,
31'b0010001010000000000000110000000,
31'b0010000000000100010000000000100,
31'b0100001000100000010000000000001,
31'b0010000000000000010000000000100,
31'b0100000000001000001010000000000,
31'b0100010000110000000000000000100,
31'b0100000000000100001010000000000,
31'b0100000000000010001010000000000,
31'b0100000000000000001010000000000,
31'b0111001000000000000010000000000,
31'b1000100001000001000000000000010,
31'b0010000000010000010000000000100,
31'b0101010000000000010000010000000,
31'b0100010000100000000000000000100,
31'b0100010000100010000000000000100,
31'b0100010000100100000000000000100,
31'b0100000000010000001010000000000,
31'b0100010000011000000000000000100,
31'b0100001000000000010000000000001,
31'b0010000000100000010000000000100,
31'b0100001000000100010000000000001,
31'b0100010000010000000000000000100,
31'b0011000000000000000000010000000,
31'b0100010000010100000000000000100,
31'b0100000000100000001010000000000,
31'b0100010000001000000000000000100,
31'b0100010000001010000000000000100,
31'b0000001000000000001000010000000,
31'b0001000000000000000010000000101,
31'b0100010000000000000000000000100,
31'b0100010000000010000000000000100,
31'b0100010000000100000000000000100,
31'b0100010000000110000000000000100,
31'b1000100000100000000010000001000,
31'b1000000000010000100000001001000,
31'b1000000010000000001000001000000,
31'b1000000000000001000010000000100,
31'b0001110000100000000001000000000,
31'b0011010000000000000000100000001,
31'b1000000010001000001000001000000,
31'b0010000010000001000100000000000,
31'b1000010000100001001000000000000,
31'b1000000000000000100000001001000,
31'b1000010000000000100010000000010,
31'b1000000000010001000010000000100,
31'b0000010000000000100000000010001,
31'b1010000000000001000000010000001,
31'b0001100100000000000000000110000,
31'b0010001000100000000000110000000,
31'b1000100000000000000010000001000,
31'b1000100000000010000010000001000,
31'b1000100000000100000010000001000,
31'b1000110000000000000000001000010,
31'b0001110000000000000001000000000,
31'b0100100001000000000000001001000,
31'b0001110000000100000001000000000,
31'b0010001000010000000000110000000,
31'b1000010000000001001000000000000,
31'b1000010000000011001000000000000,
31'b1000010000000101001000000000000,
31'b0110000000000000000101000010000,
31'b0000000000000000000000010101000,
31'b0010010000000000000100001000000,
31'b0000011100000000000000000000010,
31'b0010001000000000000000110000000,
31'b0011000000000000000001100000010,
31'b0001100000100000000000000000011,
31'b0010000010000000010000000000100,
31'b1010000000001000000000101000000,
31'b1000001000000000000000001101000,
31'b1010000000000100000000101000000,
31'b1000000000000000010110000000000,
31'b1010000000000000000000101000000,
31'b0110000100000000000001000000100,
31'b0000100100000000000000000101000,
31'b0010101100000000000000100000000,
31'b0001010000000000100000000001001,
31'b0100000000000000100010000001000,
31'b0100100000000000001000000000110,
31'b1001000000000000100000001010000,
31'b1010000000010000000000101000000,
31'b1000100001000000000010000001000,
31'b0001100000000000000000000000011,
31'b0010000010100000010000000000100,
31'b0001100000000100000000000000011,
31'b0100100000000010000000001001000,
31'b0100100000000000000000001001000,
31'b1000100000000000000001001000001,
31'b1010000000100000000000101000000,
31'b1100001100000000000000000001000,
31'b0001100000010000000000000000011,
31'b0000001010000000001000010000000,
31'b0001000000000000000000010110000,
31'b0100010010000000000000000000100,
31'b0100100000010000000000001001000,
31'b0100010010000100000000000000100,
31'b1011000000000000000100000000001,
31'b0011101000000000000000000000000,
31'b1010000000000000001100000000010,
31'b1001000000000011000001000000000,
31'b1001000000000001000001000000000,
31'b0000000000000001000000001000010,
31'b0000100000010100001000000000000,
31'b0000100000010010001000000000000,
31'b0000100000010000001000000000000,
31'b0011101000010000000000000000000,
31'b0000100000001100001000000000000,
31'b0010000100000000000001000000010,
31'b0000100000001000001000000000000,
31'b0000100000000110001000000000000,
31'b0000100000000100001000000000000,
31'b0000100000000010001000000000000,
31'b0000100000000000001000000000000,
31'b0011101000100000000000000000000,
31'b1111000000000000000000000100000,
31'b0000010010011000000000000000010,
31'b1100000001000000101000000000000,
31'b0000110000000000000010000000100,
31'b0000110000000010000010000000100,
31'b0000010010010000000000000000010,
31'b0000100000110000001000000000000,
31'b1100000011000000000000000001000,
31'b0000101000000000010010000000001,
31'b0000010010001000000000000000010,
31'b0000100000101000001000000000000,
31'b0000010010000100000000000000010,
31'b0000100000100100001000000000000,
31'b0000010010000000000000000000010,
31'b0000100000100000001000000000000,
31'b0011101001000000000000000000000,
31'b1100000000000001000010000000010,
31'b0010100010010000000000100000000,
31'b1100000000100000101000000000000,
31'b0000100000000000000000100110000,
31'b0100000000000101000000000010001,
31'b0100000000000011000000000010001,
31'b0100000000000001000000000010001,
31'b1100000010100000000000000001000,
31'b0000101010000000000000000101000,
31'b0010100010000000000000100000000,
31'b0000100001001000001000000000000,
31'b0000100001000110001000000000000,
31'b0000100001000100001000000000000,
31'b0000100001000010001000000000000,
31'b0000100001000000001000000000000,
31'b1100000010010000000000000001000,
31'b1000000000000000000101010000000,
31'b0000000100010000001000010000000,
31'b1100000000000000101000000000000,
31'b0011000000000000000010001100000,
31'b1100001000000000000000100010000,
31'b0001010100000000010010000000000,
31'b1100000000001000101000000000000,
31'b1100000010000000000000000001000,
31'b0000000010000100000001000000001,
31'b0000000100000000001000010000000,
31'b0000000010000000000001000000001,
31'b1100000010001000000000000001000,
31'b0000100001100100001000000000000,
31'b0000010011000000000000000000010,
31'b0000100001100000001000000000000,
31'b0110000000000000010000000000010,
31'b0110000000000010010000000000010,
31'b0110000000000100010000000000010,
31'b1001000010000001000001000000000,
31'b0000100000000000100000000001000,
31'b0000100000000010100000000001000,
31'b0000100000000100100000000001000,
31'b0000100010010000001000000000000,
31'b1100000001100000000000000001000,
31'b0000101001000000000000000101000,
31'b0010100001000000000000100000000,
31'b0000100010001000001000000000000,
31'b0000100000010000100000000001000,
31'b0000100010000100001000000000000,
31'b0000010000100000000000000000010,
31'b0000100010000000001000000000000,
31'b1100000001010000000000000001000,
31'b0000000101000000100000010001000,
31'b0000010000011000000000000000010,
31'b0000000001010000000001000000001,
31'b0000100000100000100000000001000,
31'b0000000000010000000010001001000,
31'b0000010000010000000000000000010,
31'b0000000000000001100000000000100,
31'b1100000001000000000000000001000,
31'b0000000001000100000001000000001,
31'b0000010000001000000000000000010,
31'b0000000001000000000001000000001,
31'b0000010000000100000000000000010,
31'b0000000000000000000010001001000,
31'b0000010000000000000000000000010,
31'b0000010000000010000000000000010,
31'b1100000000110000000000000001000,
31'b0001100000000100100000000010000,
31'b0010100000010000000000100000000,
31'b0001100000000000100000000010000,
31'b1000000000000000000100100000010,
31'b1000001000000000000010010001000,
31'b1010010000000000010000000001000,
31'b0101000000000000001001000000100,
31'b1100000000100000000000000001000,
31'b0000101000000000000000000101000,
31'b0010100000000000000000100000000,
31'b0000000000100000000001000000001,
31'b1100000000101000000000000001000,
31'b0000101000001000000000000101000,
31'b0010100000001000000000100000000,
31'b0000100011000000001000000000000,
31'b1100000000010000000000000001000,
31'b0000000100000000100000010001000,
31'b0000000000000000110100000000000,
31'b0000000000010000000001000000001,
31'b1100000000011000000000000001000,
31'b0010000100000001000000001000001,
31'b0000010001010000000000000000010,
31'b0000000001000001100000000000100,
31'b1100000000000000000000000001000,
31'b0000000000000100000001000000001,
31'b0000000000000010000001000000001,
31'b0000000000000000000001000000001,
31'b1100000000001000000000000001000,
31'b0000000001000000000010001001000,
31'b0000010001000000000000000000010,
31'b0000000000001000000001000000001,
31'b1000100000001000000101000000000,
31'b0100000010000000000010000101000,
31'b1000001000000000001000001000000,
31'b1001000100000001000001000000000,
31'b1000100000000000000101000000000,
31'b1011000000010000000000001000000,
31'b1000100000000100000101000000000,
31'b0010001000000001000100000000000,
31'b0010000000000100000001000000010,
31'b1011000000001000000000001000000,
31'b0010000000000000000001000000010,
31'b0010000000000010000001000000010,
31'b1011000000000010000000001000000,
31'b1011000000000000000000001000000,
31'b0010000000001000000001000000010,
31'b0000100100000000001000000000000,
31'b0100000001000010010000000000001,
31'b0100000001000000010000000000001,
31'b0000000001010000001000010000000,
31'b0100100000000000001000001100000,
31'b1000100000100000000101000000000,
31'b1010000000000000000100100000001,
31'b0001010001000000010010000000000,
31'b0010001000100001000100000000000,
31'b0100000000000001000000000100010,
31'b0100000001010000010000000000001,
31'b0000000001000000001000010000000,
31'b0000100000000000000000100000011,
31'b0100011001000000000000000000100,
31'b1011000000100000000000001000000,
31'b0000010110000000000000000000010,
31'b0010000010000000000000110000000,
31'b0111000000010000000010000000000,
31'b0100000000100000010000000000001,
31'b0010001000000000010000000000100,
31'b0100001000001000001010000000000,
31'b1000100001000000000101000000000,
31'b0100001000000100001010000000000,
31'b0101000000000000000000010000101,
31'b0100001000000000001010000000000,
31'b0111000000000000000010000000000,
31'b0111000000000010000010000000000,
31'b0000000000100000001000010000000,
31'b0010010000001000000000000000001,
31'b0111000000001000000010000000000,
31'b0010010000000100000000000000001,
31'b0010010000000010000000000000001,
31'b0010010000000000000000000000001,
31'b0100000000000010010000000000001,
31'b0100000000000000010000000000001,
31'b0000000000010000001000010000000,
31'b0100000000000100010000000000001,
31'b0100011000010000000000000000100,
31'b0100000000001000010000000000001,
31'b0001010000000000010010000000000,
31'b0100001000100000001010000000000,
31'b0000000000000100001000010000000,
31'b0100000000010000010000000000001,
31'b0000000000000000001000010000000,
31'b0000000000000010001000010000000,
31'b0100011000000000000000000000100,
31'b0100011000000010000000000000100,
31'b0000000000001000001000010000000,
31'b0010010000100000000000000000001,
31'b0110000100000000010000000000010,
31'b0100000000000000000010000101000,
31'b1000001010000000001000001000000,
31'b1001000000000000000000001110000,
31'b0000100100000000100000000001000,
31'b0100100000000000011001000000000,
31'b0001010000000000000000000101001,
31'b0010001010000001000100000000000,
31'b0011000000000000010000100000100,
31'b1101000000000001010000000000000,
31'b0010000010000000000001000000010,
31'b0010000010000010000001000000010,
31'b0000100100010000100000000001000,
31'b1100100000000000000000010001000,
31'b0000100000000000000001010000001,
31'b0010000000100000000000110000000,
31'b1000101000000000000010000001000,
31'b0000000001000000100000010001000,
31'b0001010000000000001100001000000,
31'b0010000000011000000000110000000,
31'b0001111000000000000001000000000,
31'b0010000001000001000000001000001,
31'b0001000000000000100000010010000,
31'b0010000000010000000000110000000,
31'b1100000101000000000000000001000,
31'b0010000000001100000000110000000,
31'b0000010100001000000000000000010,
31'b0010000000001000000000110000000,
31'b0000010100000100000000000000010,
31'b0010000000000100000000110000000,
31'b0000010100000000000000000000010,
31'b0010000000000000000000110000000,
31'b1000000000100000001100000000001,
31'b0000010000000000000000000110001,
31'b0010100100010000000000100000000,
31'b0001100100000000100000000010000,
31'b1000000000000000000000001101000,
31'b1010010000000000000100010000000,
31'b1000001000000000010110000000000,
31'b1010001000000000000000101000000,
31'b1100000100100000000000000001000,
31'b0000110000000100000000010000010,
31'b0010100100000000000000100000000,
31'b0000110000000000000000010000010,
31'b1101000000000000000100000000100,
31'b0011000000000001000100100000000,
31'b0010100100001000000000100000000,
31'b0010010010000000000000000000001,
31'b1000000000000000001100000000001,
31'b0000000000000000100000010001000,
31'b0000000100000000110100000000000,
31'b0000000100010000000001000000001,
31'b1000000000100000000000001101000,
31'b0010000000000001000000001000001,
31'b0001010010000000010010000000000,
31'b0010000001010000000000110000000,
31'b1100000100000000000000000001000,
31'b0000000100000100000001000000001,
31'b0000000010000000001000010000000,
31'b0000000100000000000001000000001,
31'b1100000100001000000000000001000,
31'b0010000001000100000000110000000,
31'b0000010101000000000000000000010,
31'b0010000001000000000000110000000,
31'b0011110000000000000000000000000,
31'b0110000010000000000100000100000,
31'b1001000001000000110000000000000,
31'b0100000010000000000010010000010,
31'b0011110000001000000000000000000,
31'b1100000000000000000010000100100,
31'b0100000000100000000011100000000,
31'b0100000000010000000100000010000,
31'b0101000001000000000100000001000,
31'b0100100000000000000000010000100,
31'b0100000000100001000000010001000,
31'b0100000000001000000100000010000,
31'b0100000101100000000000000000100,
31'b0100000000000100000100000010000,
31'b0100000000000010000100000010000,
31'b0100000000000000000100000010000,
31'b0011110000100000000000000000000,
31'b0011000010000000001000000000010,
31'b0100000000010001000000010001000,
31'b0000000010000001000101000000000,
31'b0001000001000000000000100000010,
31'b1000000001000000100000010000100,
31'b0100000000000000000011100000000,
31'b0100000000110000000100000010000,
31'b1000001000000000000000010100100,
31'b1000000100000000000010001000100,
31'b0100000000000001000000010001000,
31'b0100000000101000000100000010000,
31'b0100000101000000000000000000100,
31'b0100000101000010000000000000100,
31'b0000001010000000000000000000010,
31'b0100000000100000000100000010000,
31'b0000000000000000000000001100100,
31'b0001000010000000000001010000000,
31'b1001000000000000110000000000000,
31'b1001000000000010110000000000000,
31'b0001000000100000000000100000010,
31'b1000000010000000010000100100000,
31'b1001000000001000110000000000000,
31'b0100010100000000001010000000000,
31'b0101000000000000000100000001000,
31'b0101000000000010000100000001000,
31'b1001000000010000110000000000000,
31'b1010000000000000010000100010000,
31'b0100000100100000000000000000100,
31'b0100000100100010000000000000100,
31'b0100000100100100000000000000100,
31'b0100000001000000000100000010000,
31'b0001000000001000000000100000010,
31'b1000000000001000100000010000100,
31'b1001000000100000110000000000000,
31'b1000000000000000000001101000000,
31'b0001000000000000000000100000010,
31'b1000000000000000100000010000100,
31'b0001000000000100000000100000010,
31'b1000000000001000000001101000000,
31'b0100000100001000000000000000100,
31'b0100100000000000010000000011000,
31'b0100000100001100000000000000100,
31'b1010000000000000100010000000001,
31'b0100000100000000000000000000100,
31'b0100000100000010000000000000100,
31'b0100000100000100000000000000100,
31'b0100000100000110000000000000100,
31'b0110000000000010000100000100000,
31'b0110000000000000000100000100000,
31'b0100001000000000000100100001000,
31'b0100000000000000000010010000010,
31'b0001100100100000000001000000000,
31'b1100000000000000000000010010001,
31'b0000001000110000000000000000010,
31'b0100000010010000000100000010000,
31'b1000001000000000110000100000000,
31'b0110000000010000000100000100000,
31'b0000001000101000000000000000010,
31'b0100000010001000000100000010000,
31'b0000001000100100000000000000010,
31'b0110000000000000000000000000111,
31'b0000001000100000000000000000010,
31'b0100000010000000000100000010000,
31'b1010101000000000000100000000000,
31'b0011000000000000001000000000010,
31'b0000001000011000000000000000010,
31'b0000000000000001000101000000000,
31'b0001100100000000000001000000000,
31'b0011000000001000001000000000010,
31'b0000001000010000000000000000010,
31'b0000001000010010000000000000010,
31'b1000000100000001001000000000000,
31'b1001001000000000000001001000000,
31'b0000001000001000000000000000010,
31'b0000001000001010000000000000010,
31'b0000001000000100000000000000010,
31'b0010000100000000000100001000000,
31'b0000001000000000000000000000010,
31'b0000001000000010000000000000010,
31'b0001000000000010000001010000000,
31'b0001000000000000000001010000000,
31'b1001000010000000110000000000000,
31'b0001000000000100000001010000000,
31'b1000000000000100000000011000010,
31'b1000000000000000010000100100000,
31'b1000000000000000000000011000010,
31'b1000000000000100010000100100000,
31'b0110010000000000000001000000100,
31'b0001000000010000000001010000000,
31'b0010111000000000000000100000000,
31'b0001000100000000100000000001001,
31'b0110001000000000100100000000000,
31'b1000100000000001001000010000000,
31'b0010000000000000000000001010100,
31'b0100000100000000100000001000010,
31'b0001000010001000000000100000010,
31'b0001000000100000000001010000000,
31'b0000000000001000010001000000100,
31'b0000000000000000100000000100010,
31'b0001000010000000000000100000010,
31'b1000000010000000100000010000100,
31'b0000000000000000010001000000100,
31'b0000000000001000100000000100010,
31'b1100011000000000000000000001000,
31'b0001001000000000000000000011010,
31'b0000010000000001000000000100100,
31'b0000011000000000000001000000001,
31'b0100000110000000000000000000100,
31'b0100001000000000000000001010001,
31'b0000001001000000000000000000010,
31'b0000001001000010000000000000010,
31'b1000100000000000100000000000100,
31'b1000100000000010100000000000100,
31'b1000010000000000001000001000000,
31'b1000010000000010001000001000000,
31'b1100000000000000001001000010000,
31'b0011000010000000000000100000001,
31'b1000010000001000001000001000000,
31'b0010010000000001000100000000000,
31'b1000100000010000100000000000100,
31'b1000110000000001000000000000010,
31'b1000010000010000001000001000000,
31'b0101000001000000010000010000000,
31'b0100000001100000000000000000100,
31'b0100000100000100000100000010000,
31'b0100000100000010000100000010000,
31'b0100000100000000000100000010000,
31'b1000100000100000100000000000100,
31'b1000000000010000000010001000100,
31'b1000010000100000001000001000000,
31'b1000000000000001100000000001000,
31'b0100000001010000000000000000100,
31'b0100010000000000000101000100000,
31'b0100000100000000000011100000000,
31'b1010000000000000000000011000001,
31'b1000000010000001001000000000000,
31'b1000000000000000000010001000100,
31'b1000010000000000000000000001110,
31'b1000000000010001100000000001000,
31'b0100000001000000000000000000100,
31'b0100000001000010000000000000100,
31'b0100000001000100000000000000100,
31'b0100000100100000000100000010000,
31'b0001000000000000001000000000001,
31'b0001000000000010001000000000001,
31'b0010010000000000010000000000100,
31'b0101000000010000010000010000000,
31'b0100000000110000000000000000100,
31'b0100010000000100001010000000000,
31'b0100010000000010001010000000000,
31'b0100010000000000001010000000000,
31'b0100000000101000000000000000100,
31'b0101000000000100010000010000000,
31'b0101000000000010010000010000000,
31'b0101000000000000010000010000000,
31'b0100000000100000000000000000100,
31'b0100000000100010000000000000100,
31'b0100000000100100000000000000100,
31'b0010001000000000000000000000001,
31'b0100000000011000000000000000100,
31'b0100011000000000010000000000001,
31'b0110000000000000000010010000001,
31'b1000000100000000000001101000000,
31'b0100000000010000000000000000100,
31'b0100000000010010000000000000100,
31'b0100000000010100000000000000100,
31'b0100010000100000001010000000000,
31'b0100000000001000000000000000100,
31'b0100000000001010000000000000100,
31'b0100000000001100000000000000100,
31'b0101000000100000010000010000000,
31'b0100000000000000000000000000100,
31'b0100000000000010000000000000100,
31'b0100000000000100000000000000100,
31'b0100000000000110000000000000100,
31'b1000100010000000100000000000100,
31'b0110000100000000000100000100000,
31'b1000010010000000001000001000000,
31'b1000100000100000000000001000010,
31'b0001100000100000000001000000000,
31'b0011000000000000000000100000001,
31'b0001100000100100000001000000000,
31'b0011000000000100000000100000001,
31'b1000000000100001001000000000000,
31'b1000010000000000100000001001000,
31'b1000000000000000100010000000010,
31'b1000100000000000001000000001100,
31'b0000000000000000100000000010001,
31'b0010000000100000000100001000000,
31'b0000001100100000000000000000010,
31'b0100000110000000000100000010000,
31'b1000000000010001001000000000000,
31'b1000100000000100000000001000010,
31'b1000100000000010000000001000010,
31'b1000100000000000000000001000010,
31'b0001100000000000000001000000000,
31'b0010000000010000000100001000000,
31'b0001100000000100000001000000000,
31'b1011001000000001000000000000000,
31'b1000000000000001001000000000000,
31'b1000000000000011001000000000000,
31'b1000000000000101001000000000000,
31'b1000100000010000000000001000010,
31'b0000000000000000010010100000000,
31'b0010000000000000000100001000000,
31'b0000001100000000000000000000010,
31'b0010000000000100000100001000000,
31'b0001000010000000001000000000001,
31'b0001000100000000000001010000000,
31'b0010010010000000010000000000100,
31'b0001000100000100000001010000000,
31'b0100100000000001101000000000000,
31'b1010001000000000000100010000000,
31'b1000010000000000010110000000000,
31'b1010010000000000000000101000000,
31'b1101000000000000100001000000000,
31'b0001000100010000000001010000000,
31'b1001000000000000001100010000000,
31'b0001000000000000100000000001001,
31'b0100000010100000000000000000100,
31'b0100000010100010000000000000100,
31'b0100000010100100000000000000100,
31'b0100000000000000100000001000010,
31'b1100100000000000000000000010001,
31'b0001110000000000000000000000011,
31'b0110000000000000000000000110100,
31'b0000100000000000000001000011000,
31'b0100000010010000000000000000100,
31'b0100110000000000000000001001000,
31'b0100100000000000000010000000010,
31'b0100100000000010000010000000010,
31'b1000000001000001001000000000000,
31'b1100000000000000010000101000000,
31'b1100000000000000000000010100010,
31'b0001010000000000000000010110000,
31'b0100000010000000000000000000100,
31'b0100000010000010000000000000100,
31'b0100000010000100000000000000100,
31'b0100000010000110000000000000100,
31'b0011111000000000000000000000000,
31'b0000000101000000000010010000100,
31'b0100000010000000000100100001000,
31'b0000000000010000000001110000000,
31'b0000100000100000000010000000100,
31'b0000000000010000100000001000100,
31'b0000000010110000000000000000010,
31'b0000000000000001000010000001000,
31'b1000000010000000110000100000000,
31'b0000000000001000100000001000100,
31'b0000000010101000000000000000010,
31'b0000000000000000000001110000000,
31'b0000000010100100000000000000010,
31'b0000000000000000100000001000100,
31'b0000000010100000000000000000010,
31'b0000110000000000001000000000000,
31'b0010000000000000000000000110010,
31'b0110100000000000011000000000000,
31'b0000000010011000000000000000010,
31'b0000001010000001000101000000000,
31'b0000100000000000000010000000100,
31'b0000100000000010000010000000100,
31'b0000000010010000000000000000010,
31'b0000000010010010000000000000010,
31'b1000000000000000000000010100100,
31'b1001000010000000000001001000000,
31'b0000000010001000000000000000010,
31'b0000000010001010000000000000010,
31'b0000000010000100000000000000010,
31'b0000000010000110000000000000010,
31'b0000000010000000000000000000010,
31'b0000000010000010000000000000010,
31'b0001000000000001000010000010000,
31'b0000000100000000000010010000100,
31'b1100000000000001000000001001000,
31'b0010000100011000000000000000001,
31'b0001001000100000000000100000010,
31'b0010000100010100000000000000001,
31'b1010000010000000010000000001000,
31'b0010000100010000000000000000001,
31'b1100000000000000100010000000100,
31'b0010000100001100000000000000001,
31'b0010110010000000000000100000000,
31'b0010000100001000000000000000001,
31'b0110000010000000100100000000000,
31'b0010000100000100000000000000001,
31'b0010000100000010000000000000001,
31'b0010000100000000000000000000001,
31'b0010100000000001000000101000000,
31'b1100100000000000000000001000100,
31'b0001000100001000010010000000000,
31'b1100010000000000101000000000000,
31'b0001001000000000000000100000010,
31'b1000100000000000001100100000000,
31'b0001000100000000010010000000000,
31'b0011000000000000000000000101010,
31'b1100010010000000000000000001000,
31'b0010000000000100001000100000010,
31'b0000010100000000001000010000000,
31'b0010000000000000001000100000010,
31'b0100001100000000000000000000100,
31'b0100001100000010000000000000100,
31'b0000000011000000000000000000010,
31'b0010000100100000000000000000001,
31'b1010100000100000000100000000000,
31'b1011000000000000010000000010000,
31'b0100000000000000000100100001000,
31'b0100001000000000000010010000010,
31'b0000110000000000100000000001000,
31'b0000110000000010100000000001000,
31'b0000000000110000000000000000010,
31'b0000000010000001000010000001000,
31'b1000000000000000110000100000000,
31'b1001000000100000000001001000000,
31'b0000000000101000000000000000010,
31'b0000000010000000000001110000000,
31'b0000000000100100000000000000010,
31'b0000000010000000100000001000100,
31'b0000000000100000000000000000010,
31'b0000000000100010000000000000010,
31'b1010100000000000000100000000000,
31'b1010100000000010000100000000000,
31'b0000000000011000000000000000010,
31'b0000001000000001000101000000000,
31'b0000000000010100000000000000010,
31'b0000100000000001001000001000000,
31'b0000000000010000000000000000010,
31'b0000000000010010000000000000010,
31'b0000000000001100000000000000010,
31'b1001000000000000000001001000000,
31'b0000000000001000000000000000010,
31'b0000000000001010000000000000010,
31'b0000000000000100000000000000010,
31'b0000000000000110000000000000010,
31'b0000000000000000000000000000010,
31'b0000000000000010000000000000010,
31'b0001001000000010000001010000000,
31'b0001001000000000000001010000000,
31'b1100100000000000100000000000010,
31'b0001110000000000100000000010000,
31'b1010000000000100010000000001000,
31'b1010000100000000000100010000000,
31'b1010000000000000010000000001000,
31'b1010000000000010010000000001000,
31'b1100010000100000000000000001000,
31'b0001001000010000000001010000000,
31'b0010110000000000000000100000000,
31'b0000100100000000000000010000010,
31'b0110000000000000100100000000000,
31'b0110000000000010100100000000000,
31'b0000000001100000000000000000010,
31'b0010000110000000000000000000001,
31'b1100010000010000000000000001000,
31'b0001001000100000000001010000000,
31'b0000010000000000110100000000000,
31'b0000010000010000000001000000001,
31'b0100100000000000010000100000000,
31'b0100100000000010010000100000000,
31'b0000000001010000000000000000010,
31'b0000000001010010000000000000010,
31'b1100010000000000000000000001000,
31'b0001000000000000000000000011010,
31'b0000000001001000000000000000010,
31'b0000010000000000000001000000001,
31'b0000000001000100000000000000010,
31'b0100000000000000000000001010001,
31'b0000000001000000000000000000010,
31'b0000000001000010000000000000010,
31'b1000101000000000100000000000100,
31'b0000000001000000000010010000100,
31'b1100000000000000100001100000000,
31'b0010000001011000000000000000001,
31'b1100000000000000000000011000100,
31'b0010000001010100000000000000001,
31'b0010000001010010000000000000001,
31'b0010000001010000000000000000001,
31'b0011000000000000000000000011001,
31'b0010000001001100000000000000001,
31'b0010010000000000000001000000010,
31'b0010000001001000000000000000001,
31'b0110000000000000000000001010010,
31'b0010000001000100000000000000001,
31'b0010000001000010000000000000001,
31'b0010000001000000000000000000001,
31'b0100000000001000010001000000010,
31'b0100000000000000100000000100100,
31'b0001000010000000001100001000000,
31'b1101000000000000010000001000000,
31'b0100000000000000010001000000010,
31'b0100000000001000100000000100100,
31'b0001000001000000010010000000000,
31'b1011000010000001000000000000000,
31'b1000001010000001001000000000000,
31'b1001000000000001000000000110000,
31'b0000010001000000001000010000000,
31'b0010100010000000001001000000000,
31'b0100001001000000000000000000100,
31'b0100001001000010000000000000100,
31'b0000000110000000000000000000010,
31'b0010000001100000000000000000001,
31'b0001001000000000001000000000001,
31'b0000000000000000000010010000100,
31'b0010011000000000010000000000100,
31'b0010000000011000000000000000001,
31'b0110000000000000011000010000000,
31'b0010000000010100000000000000001,
31'b0010000000010010000000000000001,
31'b0010000000010000000000000000001,
31'b0111010000000000000010000000000,
31'b0010000000001100000000000000001,
31'b0010000000001010000000000000001,
31'b0010000000001000000000000000001,
31'b0100001000100000000000000000100,
31'b0010000000000100000000000000001,
31'b0010000000000010000000000000001,
31'b0010000000000000000000000000001,
31'b0100010000000010010000000000001,
31'b0100010000000000010000000000001,
31'b0001000000001000010010000000000,
31'b0111000000000000001000000000100,
31'b0100001000010000000000000000100,
31'b0100010000001000010000000000001,
31'b0001000000000000010010000000000,
31'b0010000000110000000000000000001,
31'b0100001000001000000000000000100,
31'b0100010000010000010000000000001,
31'b0000010000000000001000010000000,
31'b0010000000101000000000000000001,
31'b0100001000000000000000000000100,
31'b0100001000000010000000000000100,
31'b0000100000000000000001100000000,
31'b0010000000100000000000000000001,
31'b0100000000000100000000001100010,
31'b0100000000000000010000110000000,
31'b0100000000000000000000001100010,
31'b0100000000000100010000110000000,
31'b0001101000100000000001000000000,
31'b1101000000000000000001000100000,
31'b0001000000000000000000000101001,
31'b1011000000100001000000000000000,
31'b0000000000000100001000100000001,
31'b0100100000000001001000000100000,
31'b0000000000000000001000100000001,
31'b0000100001000000000000010000010,
31'b0000001000000000100000000010001,
31'b0010001000100000000100001000000,
31'b0000000100100000000000000000010,
31'b0010000011000000000000000000001,
31'b1010100100000000000100000000000,
31'b0100000010000000100000000100100,
31'b0001000000000000001100001000000,
31'b1011000000001001000000000000000,
31'b0001101000000000000001000000000,
31'b1011000000000101000000000000000,
31'b0000000100010000000000000000010,
31'b1011000000000001000000000000000,
31'b1000001000000001001000000000000,
31'b1001000100000000000001001000000,
31'b0000000100001000000000000000010,
31'b0010100000000000001001000000000,
31'b0000000100000100000000000000010,
31'b0010001000000000000100001000000,
31'b0000000100000000000000000000010,
31'b0000000100000010000000000000010,
31'b0000000000000010000000000110001,
31'b0000000000000000000000000110001,
31'b0100100000000001000000100010000,
31'b0000100000010000000000010000010,
31'b1010000000000010000100010000000,
31'b1010000000000000000100010000000,
31'b1010000100000000010000000001000,
31'b1000000000000000000010000100010,
31'b0000100000000110000000010000010,
31'b0000100000000100000000010000010,
31'b0000100000000010000000010000010,
31'b0000100000000000000000010000010,
31'b0110000100000000100100000000000,
31'b0010000010000100000000000000001,
31'b0010000010000010000000000000001,
31'b0010000010000000000000000000001,
31'b1010000000000001000000000011000,
31'b0000010000000000100000010001000,
31'b0001000010001000010010000000000,
31'b0000101000000000000001000011000,
31'b0100100100000000010000100000000,
31'b1010000000100000000100010000000,
31'b0001000010000000010010000000000,
31'b1011000001000001000000000000000,
31'b1100010100000000000000000001000,
31'b0001100000000000100001000100000,
31'b0000010010000000001000010000000,
31'b0000100000100000000000010000010,
31'b0100001010000000000000000000100,
31'b0100001010000010000000000000100,
31'b0000000101000000000000000000010,
31'b0010000010100000000000000000001,
31'b0100000000000000000000000000000,
31'b0100000000000010000000000000000,
31'b0100000000000100000000000000000,
31'b0100000000000110000000000000000,
31'b0100000000001000000000000000000,
31'b0100000000001010000000000000000,
31'b0100000000001100000000000000000,
31'b0100000000001110000000000000000,
31'b0100000000010000000000000000000,
31'b0100000000010010000000000000000,
31'b0100000000010100000000000000000,
31'b0100000000010110000000000000000,
31'b0100000000011000000000000000000,
31'b0100000000011010000000000000000,
31'b0100000000011100000000000000000,
31'b0111001000000000001000000000000,
31'b0100000000100000000000000000000,
31'b0100000000100010000000000000000,
31'b0100000000100100000000000000000,
31'b0100000000100110000000000000000,
31'b0100000000101000000000000000000,
31'b0100000000101010000000000000000,
31'b0100000000101100000000000000000,
31'b0101000000000000010000010000100,
31'b0100000000110000000000000000000,
31'b0100000000110010000000000000000,
31'b0100000000110100000000000000000,
31'b0100010000000000001010000000100,
31'b0000000100000000000000001100000,
31'b0000001000000000000010010000000,
31'b0010010000000000010000000000000,
31'b0010010000000010010000000000000,
31'b0100000001000000000000000000000,
31'b0100000001000010000000000000000,
31'b0100000001000100000000000000000,
31'b0100000001000110000000000000000,
31'b0100000001001000000000000000000,
31'b1000000000000000000010001000000,
31'b1000010000000000000000000001010,
31'b1000000000000100000010001000000,
31'b0100000001010000000000000000000,
31'b0100000001010010000000000000000,
31'b0100000001010100000000000000000,
31'b0100000001010110000000000000000,
31'b1000100000100000100000000000000,
31'b1000000000010000000010001000000,
31'b1000100000100100100000000000000,
31'b1000000000010100000010001000000,
31'b0100000001100000000000000000000,
31'b0100000001100010000000000000000,
31'b0100000001100100000000000000000,
31'b0100000100000000000100000010100,
31'b1000100000010000100000000000000,
31'b1000000000100000000010001000000,
31'b1000100000010100100000000000000,
31'b1000100010000000001000000001000,
31'b1000100000001000100000000000000,
31'b1100000100000000000010000100000,
31'b1100010000000000000100100000000,
31'b0010010000000001000100000000100,
31'b1000100000000000100000000000000,
31'b1000100000000010100000000000000,
31'b1000100000000100100000000000000,
31'b1000100000000110100000000000000,
31'b0100000010000000000000000000000,
31'b0100000010000010000000000000000,
31'b0100000010000100000000000000000,
31'b0100000010000110000000000000000,
31'b0100000010001000000000000000000,
31'b0100000010001010000000000000000,
31'b0100000010001100000000000000000,
31'b0101000000000000100000100100000,
31'b0100000010010000000000000000000,
31'b0100000010010010000000000000000,
31'b0000000100000000010001000000000,
31'b0100000000000000101000000001000,
31'b0100000010011000000000000000000,
31'b0100001000000000000000100011000,
31'b0110000000000000000000000110000,
31'b0110000000000010000000000110000,
31'b0100000010100000000000000000000,
31'b0100000010100010000000000000000,
31'b0100000010100100000000000000000,
31'b0100000010100110000000000000000,
31'b0100000010101000000000000000000,
31'b0100000010101010000000000000000,
31'b0100000010101100000000000000000,
31'b1000100001000000001000000001000,
31'b0100000010110000000000000000000,
31'b0100000010110010000000000000000,
31'b0100010000000001000000001000000,
31'b0100010000000011000000001000000,
31'b0000000000000001000001000010000,
31'b0000001010000000000010010000000,
31'b0010010010000000010000000000000,
31'b1010101000000000000000000010000,
31'b0100000011000000000000000000000,
31'b0100000011000010000000000000000,
31'b0100000011000100000000000000000,
31'b0110001000000000100000000010000,
31'b1000000000000001001000000000100,
31'b1000000010000000000010001000000,
31'b1000010010000000000000000001010,
31'b1000100000100000001000000001000,
31'b0100000011010000000000000000000,
31'b0111000000000000000000000101000,
31'b0101001000000000000000100000000,
31'b0101001000000010000000100000000,
31'b1000100010100000100000000000000,
31'b1000010000000000101000000000010,
31'b0110000001000000000000000110000,
31'b1000100000000000000000001000110,
31'b0100000011100000000000000000000,
31'b0110000100000000000000000000011,
31'b0100001000000000000100001000001,
31'b1000100000001000001000000001000,
31'b1000100010010000100000000000000,
31'b1000100000000100001000000001000,
31'b1000100000000010001000000001000,
31'b1000100000000000001000000001000,
31'b1101000000000001000000000000001,
31'b0011000000000000000000100000101,
31'b0101001000100000000000100000000,
31'b0001000000000001000001000001000,
31'b1000100010000000100000000000000,
31'b1000100010000010100000000000000,
31'b1000100010000100100000000000000,
31'b1000010000000001000010000000000,
31'b0100000100000000000000000000000,
31'b0100000100000010000000000000000,
31'b0100000100000100000000000000000,
31'b0100000100000110000000000000000,
31'b0100000100001000000000000000000,
31'b0100000100001010000000000000000,
31'b0100000100001100000000000000000,
31'b0101100000000001000100000000000,
31'b0100000100010000000000000000000,
31'b1000000000000000100000010000000,
31'b0000000010000000010001000000000,
31'b1000000000000100100000010000000,
31'b0000000000100000000000001100000,
31'b1000000000001000100000010000000,
31'b0000000010001000010001000000000,
31'b1000000000001100100000010000000,
31'b0100000100100000000000000000000,
31'b0100000100100010000000000000000,
31'b0100000100100100000000000000000,
31'b0100000100100110000000000000000,
31'b0000000000010000000000001100000,
31'b0100100001000000000000010000000,
31'b0100000000000001010000000010000,
31'b0100100001000100000000010000000,
31'b0000000000001000000000001100000,
31'b1000000000100000100000010000000,
31'b0000000010100000010001000000000,
31'b1001000000000000000001000100010,
31'b0000000000000000000000001100000,
31'b0000000000000010000000001100000,
31'b0000000000000100000000001100000,
31'b0000000000000110000000001100000,
31'b0100000101000000000000000000000,
31'b0100000101000010000000000000000,
31'b0100000101000100000000000000000,
31'b0100000101000110000000000000000,
31'b1000001000000000000000010100000,
31'b1000000100000000000010001000000,
31'b1000010100000000000000000001010,
31'b1010000000000000000000110001000,
31'b0000101000000000000010000000000,
31'b1000000001000000100000010000000,
31'b0000101000000100000010000000000,
31'b1010000000000001000011000000000,
31'b0000101000001000000010000000000,
31'b1000000100010000000010001000000,
31'b0000101000001100000010000000000,
31'b0011010000000001000000000001000,
31'b0100000101100000000000000000000,
31'b0000001000000000100000001000000,
31'b0100000101100100000000000000000,
31'b0100000000000000000100000010100,
31'b0100100000000010000000010000000,
31'b0100100000000000000000010000000,
31'b0100100000000110000000010000000,
31'b0100100000000100000000010000000,
31'b0000101000100000000010000000000,
31'b1100000000000000000010000100000,
31'b0000101000100100000010000000000,
31'b1100000000000100000010000100000,
31'b0000000001000000000000001100000,
31'b0100100000010000000000010000000,
31'b0000100000000000011000000000001,
31'b0100100000010100000000010000000,
31'b0100000110000000000000000000000,
31'b0100000110000010000000000000000,
31'b0000000000010000010001000000000,
31'b0000000000000000100100000000001,
31'b0100000110001000000000000000000,
31'b0100110000000000000000100000001,
31'b0000010000000001000000000100000,
31'b0000010000000011000000000100000,
31'b0000000000000100010001000000000,
31'b1000000010000000100000010000000,
31'b0000000000000000010001000000000,
31'b0000000000000010010001000000000,
31'b0000000010100000000000001100000,
31'b1001000000000000010000001000010,
31'b0000000000001000010001000000000,
31'b0000000000001010010001000000000,
31'b0100000110100000000000000000000,
31'b0110000001000000000000000000011,
31'b0010000000000000000000001010000,
31'b0010000000000010000000001010000,
31'b0110010000000000000001000000000,
31'b0110010000000010000001000000000,
31'b0010000000001000000000001010000,
31'b1010010000000000000000000001001,
31'b0000000010001000000000001100000,
31'b1000000010100000100000010000000,
31'b0000000000100000010001000000000,
31'b0001000000000000100000101000000,
31'b0000000010000000000000001100000,
31'b0001000000000000000001010000100,
31'b0000000010000100000000001100000,
31'b0001000000001000100000101000000,
31'b0100000111000000000000000000000,
31'b0110000000100000000000000000011,
31'b0000001000000000000000000000110,
31'b0000001000000010000000000000110,
31'b1000001010000000000000010100000,
31'b1001000000000000001000010010000,
31'b0000010001000001000000000100000,
31'b0000010001000011000000000100000,
31'b0000101010000000000010000000000,
31'b1000010000000000010010000010000,
31'b0000000001000000010001000000000,
31'b0000011000000001100000000000000,
31'b0000101010001000000010000000000,
31'b0011000000000000001000000000110,
31'b0000001000000000000100000100001,
31'b0000010000000000010000000000011,
31'b0110000000000010000000000000011,
31'b0110000000000000000000000000011,
31'b0010000001000000000000001010000,
31'b0110000000000100000000000000011,
31'b0110010001000000000001000000000,
31'b0100100010000000000000010000000,
31'b0011010000000000000010000000010,
31'b1110000000000000000010000010000,
31'b0000101010100000000010000000000,
31'b1100000010000000000010000100000,
31'b0000001000000000001000001001000,
31'b0001000100000001000001000001000,
31'b0000100000000000000101000001000,
31'b0110000000000000000100000100100,
31'b0000100010000000011000000000001,
31'b1100100000000000000100000000001,
31'b0100001000000000000000000000000,
31'b0100001000000010000000000000000,
31'b0100001000000100000000000000000,
31'b0100001000000110000000000000000,
31'b0100001000001000000000000000000,
31'b0100001000001010000000000000000,
31'b0100001000001100000000000000000,
31'b0111000000010000001000000000000,
31'b0100001000010000000000000000000,
31'b0100001000010010000000000000000,
31'b0100001000010100000000000000000,
31'b0111000000001000001000000000000,
31'b0100001000011000000000000000000,
31'b0000000000100000000010010000000,
31'b0111000000000010001000000000000,
31'b0111000000000000001000000000000,
31'b0100001000100000000000000000000,
31'b1000100000000000000000000100000,
31'b0100001000100100000000000000000,
31'b0010000000000000000000000000101,
31'b0100001000101000000000000000000,
31'b0000000000010000000010010000000,
31'b0100001000101100000000000000000,
31'b0010000000001000000000000000101,
31'b0100001000110000000000000000000,
31'b0000000000001000000010010000000,
31'b0101010000000000000000010000001,
31'b0010000000010000000000000000101,
31'b0000000000000010000010010000000,
31'b0000000000000000000010010000000,
31'b0010011000000000010000000000000,
31'b0000000000000100000010010000000,
31'b0100001001000000000000000000000,
31'b0100001001000010000000000000000,
31'b0100001001000100000000000000000,
31'b0110000010000000100000000010000,
31'b1000000100000000000000010100000,
31'b1000001000000000000010001000000,
31'b1000011000000000000000000001010,
31'b1000001000000100000010001000000,
31'b0000100100000000000010000000000,
31'b0100000000001000100000000100000,
31'b0101000010000000000000100000000,
31'b0101000010000010000000100000000,
31'b0100000000000010100000000100000,
31'b0100000000000000100000000100000,
31'b0101000010001000000000100000000,
31'b0100000000000100100000000100000,
31'b0100001001100000000000000000000,
31'b0000000100000000100000001000000,
31'b0100001001100100000000000000000,
31'b0010000001000000000000000000101,
31'b1000101000010000100000000000000,
31'b0000000100001000100000001000000,
31'b0010010000000000000001000000110,
31'b0010000001001000000000000000101,
31'b1100000000000000000000011000000,
31'b0000000100010000100000001000000,
31'b1100000000000100000000011000000,
31'b0010000001010000000000000000101,
31'b1000101000000000100000000000000,
31'b0000000001000000000010010000000,
31'b1000101000000100100000000000000,
31'b0010000000000001100001000000000,
31'b0100001010000000000000000000000,
31'b0100001010000010000000000000000,
31'b0100001010000100000000000000000,
31'b0110000001000000100000000010000,
31'b0100001010001000000000000000000,
31'b0100001010001010000000000000000,
31'b0100001010001100000000000000000,
31'b1000100000000000010001001000000,
31'b0100001010010000000000000000000,
31'b0100001010010010000000000000000,
31'b0101000001000000000000100000000,
31'b0101000001000010000000100000000,
31'b0100001010011000000000000000000,
31'b0100000000000000000000100011000,
31'b1011000000000000010100000000000,
31'b1010100000100000000000000010000,
31'b0100001010100000000000000000000,
31'b0000000000000000000100000010010,
31'b0100001010100100000000000000000,
31'b0010000010000000000000000000101,
31'b0100001010101000000000000000000,
31'b0000000010010000000010010000000,
31'b1001100000000000100000100000000,
31'b1000000000000000000110000000001,
31'b0100001010110000000000000000000,
31'b0000000010001000000010010000000,
31'b0101000001100000000000100000000,
31'b1010100000001000000000000010000,
31'b0000001000000001000001000010000,
31'b0000000010000000000010010000000,
31'b1010100000000010000000000010000,
31'b1010100000000000000000000010000,
31'b0100001011000000000000000000000,
31'b0110000000000100100000000010000,
31'b0000000100000000000000000000110,
31'b0110000000000000100000000010000,
31'b1000001000000001001000000000100,
31'b1000001010000000000010001000000,
31'b0100000000000000001000000101000,
31'b0110000000001000100000000010000,
31'b0101000000000100000000100000000,
31'b0101000000000110000000100000000,
31'b0101000000000000000000100000000,
31'b0101000000000010000000100000000,
31'b0101000000001100000000100000000,
31'b0100000010000000100000000100000,
31'b0101000000001000000000100000000,
31'b0101000000001010000000100000000,
31'b0100001011100000000000000000000,
31'b0000000110000000100000001000000,
31'b0100000000000000000100001000001,
31'b0110000000100000100000000010000,
31'b0011010000000000010000100000000,
31'b0001010000000000000110001000000,
31'b0001000000000000000100000001010,
31'b1000101000000000001000000001000,
31'b1100000010000000000000011000000,
31'b0000010100000000001010000000010,
31'b0101000000100000000000100000000,
31'b0101000000100010000000100000000,
31'b1010000000000001010000010000000,
31'b0000010000000000110000000010000,
31'b0101000000101000000000100000000,
31'b1010100001000000000000000010000,
31'b0100001100000000000000000000000,
31'b0100001100000010000000000000000,
31'b0100001100000100000000000000000,
31'b0110000000000000000100001000010,
31'b1000000001000000000000010100000,
31'b1100100000010000000000001000000,
31'b1100000000000001001000000000010,
31'b0011000000000000000100000001001,
31'b0000100001000000000010000000000,
31'b1000001000000000100000010000000,
31'b0000100001000100000010000000000,
31'b1000110000000000000001000010000,
31'b0000100001001000000010000000000,
31'b1100100000000000000000001000000,
31'b0000100001001100000010000000000,
31'b1100100000000100000000001000000,
31'b0100001100100000000000000000000,
31'b0000000001000000100000001000000,
31'b0100001100100100000000000000000,
31'b0010000100000000000000000000101,
31'b1100000000000000100010000000000,
31'b0000000100010000000010010000000,
31'b1100000000000100100010000000000,
31'b0010000100001000000000000000101,
31'b0000100001100000000010000000000,
31'b0000000100001000000010010000000,
31'b0000100001100100000010000000000,
31'b0010000100010000000000000000101,
31'b0000001000000000000000001100000,
31'b0000000100000000000010010000000,
31'b0000001000000100000000001100000,
31'b0010000000000000000000101001000,
31'b0000100000010000000010000000000,
31'b0000000000100000100000001000000,
31'b0000000010000000000000000000110,
31'b0000000010000010000000000000110,
31'b1000000000000000000000010100000,
31'b1000000000000010000000010100000,
31'b1000000000000100000000010100000,
31'b1000000000000110000000010100000,
31'b0000100000000000000010000000000,
31'b0000100000000010000010000000000,
31'b0000100000000100000010000000000,
31'b0000100000000110000010000000000,
31'b0000100000001000000010000000000,
31'b0100000100000000100000000100000,
31'b0000100000001100000010000000000,
31'b0101110000000000000000000000001,
31'b0000000000000010100000001000000,
31'b0000000000000000100000001000000,
31'b0000000010100000000000000000110,
31'b0000000000000100100000001000000,
31'b1000000000100000000000010100000,
31'b0000000000001000100000001000000,
31'b1001000000000000100001000000010,
31'b0000000000001100100000001000000,
31'b0000100000100000000010000000000,
31'b0000000000010000100000001000000,
31'b0000100000100100000010000000000,
31'b0000000000010100100000001000000,
31'b0000100000101000000010000000000,
31'b0000000101000000000010010000000,
31'b0000101000000000011000000000001,
31'b0010000100000001100001000000000,
31'b0100001110000000000000000000000,
31'b0100001110000010000000000000000,
31'b0000000001000000000000000000110,
31'b0000001000000000100100000000001,
31'b1100010000000000000000000001100,
31'b0011000000000000011001000000000,
31'b0000011000000001000000000100000,
31'b0000010000000000000001000000101,
31'b0000100011000000000010000000000,
31'b1010100000000001010000000000000,
31'b0000001000000000010001000000000,
31'b0000010001000001100000000000000,
31'b0000100011001000000010000000000,
31'b1100100010000000000000001000000,
31'b0000001000001000010001000000000,
31'b0000010001001001100000000000000,
31'b0110000000000000100100000000100,
31'b0000000100000000000100000010010,
31'b0010001000000000000000001010000,
31'b0010001000000010000000001010000,
31'b1100000010000000100010000000000,
31'b0001000001000000010000010000010,
31'b0010110000000000000000100000100,
31'b1100110000000001000000000000000,
31'b0000100011100000000010000000000,
31'b0001010000000000100100010000000,
31'b0000001000100000010001000000000,
31'b0101010000000000001001000000000,
31'b0000001010000000000000001100000,
31'b0001000000000000001000001010000,
31'b0000001010000100000000001100000,
31'b1100000000000000001010000001000,
31'b0000000000000100000000000000110,
31'b0000000010100000100000001000000,
31'b0000000000000000000000000000110,
31'b0000000000000010000000000000110,
31'b1000000010000000000000010100000,
31'b1001000000000000000001001000100,
31'b0000000000001000000000000000110,
31'b0000000000001010000000000000110,
31'b0000100010000000000010000000000,
31'b0000100010000010000010000000000,
31'b0000000000010000000000000000110,
31'b0000010000000001100000000000000,
31'b0000100010001000000010000000000,
31'b0100100000000001000100100000000,
31'b0000000000000000000100000100001,
31'b0000010000001001100000000000000,
31'b0000000010000010100000001000000,
31'b0000000010000000100000001000000,
31'b0000000000100000000000000000110,
31'b0000000010000100100000001000000,
31'b1000000010100000000000010100000,
31'b0001000000000000010000010000010,
31'b0001000000000000000000101100000,
31'b0001000000000100010000010000010,
31'b0000100010100000000010000000000,
31'b0000010000000000001010000000010,
31'b0000000000000000001000001001000,
31'b0000010000100001100000000000000,
31'b0000101000000000000101000001000,
31'b0001000001000000001000001010000,
31'b0000000000100000000100000100001,
31'b1010000000000001000100000001000,
31'b0100010000000000000000000000000,
31'b0100010000000010000000000000000,
31'b0100010000000100000000000000000,
31'b0100010000000110000000000000000,
31'b0100010000001000000000000000000,
31'b0100010000001010000000000000000,
31'b0000000000000000000001001010000,
31'b0001000000000000000010000000001,
31'b0100010000010000000000000000000,
31'b0100010000010010000000000000000,
31'b0100010000010100000000000000000,
31'b0100010000010110000000000000000,
31'b0100010000011000000000000000000,
31'b0100010000011010000000000000000,
31'b0010000000100000010000000000000,
31'b0010000000100010010000000000000,
31'b0100010000100000000000000000000,
31'b0100010000100010000000000000000,
31'b0100010000100100000000000000000,
31'b0100010000100110000000000000000,
31'b0100010000101000000000000000000,
31'b0110000000000000001000010000001,
31'b0010000000010000010000000000000,
31'b0010000000010010010000000000000,
31'b0100010000110000000000000000000,
31'b0100010000110010000000000000000,
31'b0010000000001000010000000000000,
31'b0100000000000000001010000000100,
31'b0010000000000100010000000000000,
31'b0010000000000110010000000000000,
31'b0010000000000000010000000000000,
31'b0010000000000010010000000000000,
31'b0100010001000000000000000000000,
31'b0100010001000010000000000000000,
31'b1000000000001000000000000001010,
31'b1100000000000000000011000010000,
31'b1000000000000100000000000001010,
31'b1000010000000000000010001000000,
31'b1000000000000000000000000001010,
31'b1000000000000010000000000001010,
31'b0100010001010000000000000000000,
31'b0100010001010010000000000000000,
31'b1100000000100000000100100000000,
31'b0010100100000000010000010000000,
31'b1000110000100000100000000000000,
31'b1000010000010000000010001000000,
31'b1000000000010000000000000001010,
31'b1000000010100001000010000000000,
31'b0100010001100000000000000000000,
31'b0100010001100010000000000000000,
31'b1100000000010000000100100000000,
31'b0010001000000000110000000100000,
31'b1000110000010000100000000000000,
31'b1000100000000001000000000000110,
31'b1000000000100000000000000001010,
31'b1000000010010001000010000000000,
31'b1100000000000100000100100000000,
31'b0011000000000000010000000011000,
31'b1100000000000000000100100000000,
31'b0010000000000001000100000000100,
31'b1000110000000000100000000000000,
31'b1000110000000010100000000000000,
31'b0010000001000000010000000000000,
31'b1000000010000001000010000000000,
31'b0100010010000000000000000000000,
31'b0100010010000010000000000000000,
31'b0100010010000100000000000000000,
31'b0100100000000001100010000000000,
31'b0100010010001000000000000000000,
31'b0100100100000000000000100000001,
31'b0000000100000001000000000100000,
31'b0001000010000000000010000000001,
31'b0100010010010000000000000000000,
31'b0100100000000000000000001001100,
31'b0100000000100001000000001000000,
31'b0100010000000000101000000001000,
31'b0100010010011000000000000000000,
31'b1001000000000000000110010000000,
31'b0010000010100000010000000000000,
31'b1011000000000000000000000100010,
31'b0000000000000000010000000110000,
31'b0100100000000000001000000000010,
31'b0100000000010001000000001000000,
31'b0100100000000100001000000000010,
31'b0110000100000000000001000000000,
31'b0110000100000010000001000000000,
31'b0010000010010000010000000000000,
31'b1010000100000000000000000001001,
31'b0100000000000101000000001000000,
31'b0100100000010000001000000000010,
31'b0100000000000001000000001000000,
31'b0100000000000011000000001000000,
31'b0010000010000100010000000000000,
31'b1010000000000000100001010000000,
31'b0010000010000000010000000000000,
31'b1000000001000001000010000000000,
31'b0100010011000000000000000000000,
31'b0110100000000000000001010000000,
31'b1100001000000001000000010000000,
31'b0010100000000000101100000000000,
31'b1000010000000001001000000000100,
31'b1000010010000000000010001000000,
31'b1000000010000000000000000001010,
31'b1000000010000010000000000001010,
31'b0101000000000000000100011000000,
31'b1000000100000000010010000010000,
31'b0101011000000000000000100000000,
31'b0000001100000001100000000000000,
31'b1000100000000000000010000001100,
31'b1000000000000000101000000000010,
31'b1000000010010000000000000001010,
31'b1000000000100001000010000000000,
31'b0100000000000000000000110000001,
31'b0100100001000000001000000000010,
31'b0100000001010001000000001000000,
31'b0000100000000001000000010100000,
31'b0110000101000000000001000000000,
31'b1000000000010101000010000000000,
31'b1000000010100000000000000001010,
31'b1000000000010001000010000000000,
31'b0100000001000101000000001000000,
31'b0000000000000100011000100000000,
31'b0100000001000001000000001000000,
31'b0000000000000000011000100000000,
31'b1000110010000000100000000000000,
31'b1000000000000101000010000000000,
31'b1000000000000011000010000000000,
31'b1000000000000001000010000000000,
31'b0100010100000000000000000000000,
31'b0100010100000010000000000000000,
31'b0100010100000100000000000000000,
31'b0100010100000110000000000000000,
31'b0100010100001000000000000000000,
31'b0100100010000000000000100000001,
31'b0000000010000001000000000100000,
31'b0001000100000000000010000000001,
31'b0010000000000001000000000010000,
31'b1000010000000000100000010000000,
31'b0010000000000101000000000010000,
31'b1000101000000000000001000010000,
31'b0010000000001001000000000010000,
31'b1000010000001000100000010000000,
31'b0010000100100000010000000000000,
31'b0011000001000001000000000001000,
31'b0100010100100000000000000000000,
31'b0100010100100010000000000000000,
31'b0100010100100100000000000000000,
31'b1001001000000000100000000000001,
31'b0110000010000000000001000000000,
31'b0110000010000010000001000000000,
31'b0010000100010000010000000000000,
31'b1010000010000000000000000001001,
31'b0010000000100001000000000010000,
31'b1000010000100000100000010000000,
31'b0100000000000000000001000110000,
31'b0100000100000000001010000000100,
31'b0000010000000000000000001100000,
31'b0010000000000000000100010001000,
31'b0010000100000000010000000000000,
31'b0010000100000010010000000000000,
31'b0100010101000000000000000000000,
31'b0100010101000010000000000000000,
31'b1100000000000000001000000100100,
31'b0010100000010000010000010000000,
31'b1000011000000000000000010100000,
31'b1000010100000000000010001000000,
31'b1000000100000000000000000001010,
31'b1010000000000000010010000100000,
31'b0010000001000001000000000010000,
31'b1000010001000000100000010000000,
31'b0010100000000010010000010000000,
31'b0010100000000000010000010000000,
31'b0011100000100000000000000000100,
31'b0011000000000101000000000001000,
31'b1001000000100000000000000100001,
31'b0011000000000001000000000001000,
31'b0100010101100000000000000000000,
31'b0100000000000000001001100000000,
31'b1001000000000000000100000000110,
31'b0000101000000000001000000000100,
31'b0110000011000000000001000000000,
31'b0100110000000000000000010000000,
31'b1001000000010000000000000100001,
31'b0100110000000100000000010000000,
31'b0011100000001000000000000000100,
31'b1100010000000000000010000100000,
31'b1100000100000000000100100000000,
31'b0010100000100000010000010000000,
31'b0011100000000000000000000000100,
31'b0101000000000000000001000101000,
31'b1001000000000000000000000100001,
31'b1001000000000010000000000100001,
31'b0100010110000000000000000000000,
31'b0100100000001000000000100000001,
31'b0000000000001001000000000100000,
31'b0000010000000000100100000000001,
31'b0000000000000101000000000100000,
31'b0100100000000000000000100000001,
31'b0000000000000001000000000100000,
31'b0000000000000011000000000100000,
31'b0010000010000001000000000010000,
31'b1000010010000000100000010000000,
31'b0000010000000000010001000000000,
31'b0000010000000010010001000000000,
31'b0100000000000000010000001010000,
31'b0100100000010000000000100000001,
31'b0000000000010001000000000100000,
31'b0000000001000000010000000000011,
31'b0110000000001000000001000000000,
31'b0110000000001010000001000000000,
31'b0010010000000000000000001010000,
31'b1010000000001000000000000001001,
31'b0110000000000000000001000000000,
31'b0110000000000010000001000000000,
31'b0000000000100001000000000100000,
31'b1010000000000000000000000001001,
31'b0110000000011000000001000000000,
31'b1000000001000000100000100000001,
31'b0100000100000001000000001000000,
31'b0101001000000000001001000000000,
31'b0110000000010000000001000000000,
31'b0110000000010010000001000000000,
31'b0010000110000000010000000000000,
31'b1010000000010000000000000001001,
31'b0100010111000000000000000000000,
31'b1001000000000000100100001000000,
31'b0000011000000000000000000000110,
31'b0000001000010001100000000000000,
31'b0100000000000000001000010000010,
31'b0100100001000000000000100000001,
31'b0000000001000001000000000100000,
31'b0000000001000011000000000100000,
31'b1010100000000000100001000000000,
31'b1000000000000000010010000010000,
31'b0000010001000000010001000000000,
31'b0000001000000001100000000000000,
31'b0100000001000000010000001010000,
31'b0000000000000100010000000000011,
31'b0000000001010001000000000100000,
31'b0000000000000000010000000000011,
31'b1011000000000000000000000010001,
31'b1010000000000000000011001000000,
31'b0011000000001000000010000000010,
31'b0000101010000000001000000000100,
31'b0110000001000000000001000000000,
31'b0110000001000010000001000000000,
31'b0011000000000000000010000000010,
31'b1010000001000000000000000001001,
31'b1001100000000000000110000000000,
31'b1000000000000000100000100000001,
31'b0100000101000001000000001000000,
31'b0000001000100001100000000000000,
31'b0110000001010000000001000000000,
31'b1000000100000101000010000000000,
31'b1001000010000000000000000100001,
31'b1000000100000001000010000000000,
31'b0100011000000000000000000000000,
31'b0100011000000010000000000000000,
31'b0100011000000100000000000000000,
31'b0110000000000000010010010000000,
31'b0100011000001000000000000000000,
31'b0100011000001010000000000000000,
31'b0000000000000000001000010000100,
31'b0001001000000000000010000000001,
31'b0100011000010000000000000000000,
31'b0100011000010010000000000000000,
31'b0101000000100000000000010000001,
31'b1000100100000000000001000010000,
31'b0100011000011000000000000000000,
31'b0100000000000000010000000000101,
31'b0010001000100000010000000000000,
31'b0111010000000000001000000000000,
31'b0100011000100000000000000000000,
31'b0001000000000000011000000000000,
31'b0101000000010000000000010000001,
31'b0010010000000000000000000000101,
31'b0111000000000000000010000000100,
31'b0001000000001000011000000000000,
31'b0010001000010000010000000000000,
31'b0010010000001000000000000000101,
31'b0101000000000100000000010000001,
31'b0001000000010000011000000000000,
31'b0101000000000000000000010000001,
31'b0101000000000010000000010000001,
31'b0010001000000100010000000000000,
31'b0000010000000000000010010000000,
31'b0010001000000000010000000000000,
31'b0010001000000010010000000000000,
31'b0100011001000000000000000000000,
31'b0100011001000010000000000000000,
31'b1100000010000001000000010000000,
31'b0010000010000000000000110000100,
31'b1000010100000000000000010100000,
31'b1010000000000000000000100100010,
31'b1000001000000000000000000001010,
31'b1000001000000010000000000001010,
31'b0100000000000001000100000000001,
31'b0100010000001000100000000100000,
31'b0101010010000000000000100000000,
31'b0000100000000000000100100100000,
31'b0100010000000010100000000100000,
31'b0100010000000000100000000100000,
31'b1000001000010000000000000001010,
31'b0101100100000000000000000000001,
31'b0101000000000001000000101000000,
31'b0001000001000000011000000000000,
31'b0010000000001000000001000000110,
31'b0010000000000000110000000100000,
31'b0011000010000000010000100000000,
31'b0001000010000000000110001000000,
31'b0010000000000000000001000000110,
31'b0100100000000000000000000101010,
31'b1100010000000000000000011000000,
31'b0001000001010000011000000000000,
31'b1100001000000000000100100000000,
31'b0010001000000001000100000000100,
31'b1000111000000000100000000000000,
31'b0000010001000000000010010000000,
31'b1000000000000000000001010010000,
31'b1000001010000001000010000000000,
31'b1000000000000000001000000100010,
31'b1100100000000000010000000010000,
31'b1100000001000001000000010000000,
31'b0010000001000000000000110000100,
31'b1100000100000000000000000001100,
31'b0010000100000001000000100001000,
31'b0000001100000001000000000100000,
31'b0000000100000000000001000000101,
31'b1100000000000000000000101000001,
31'b0010000100000000000011010000000,
31'b0101010001000000000000100000000,
31'b0000000101000001100000000000000,
31'b1001000000000000000000100001010,
31'b0000000001000000000010100000001,
31'b0010100000000000001100000100000,
31'b0000000101001001100000000000000,
31'b1101000000000000000100000000000,
31'b0001000010000000011000000000000,
31'b1101000000000100000100000000000,
31'b0010010010000000000000000000101,
31'b1101000000001000000100000000000,
31'b0001000010001000011000000000000,
31'b0010100100000000000000100000100,
31'b1100100100000001000000000000000,
31'b1101000000010000000100000000000,
31'b0001000100000000100100010000000,
31'b0100001000000001000000001000000,
31'b0101000100000000001001000000000,
31'b0010100001000000000011000000000,
31'b0000010010000000000010010000000,
31'b0010001010000000010000000000000,
31'b1010110000000000000000000010000,
31'b1100000000000101000000010000000,
31'b0010000000001000100001001000000,
31'b1100000000000001000000010000000,
31'b0010000000000000000000110000100,
31'b0011000000100000010000100000000,
31'b0010000000000000100001001000000,
31'b1100000000001001000000010000000,
31'b0010000000001000000000110000100,
31'b0101010000000100000000100000000,
31'b0000000100000101100000000000000,
31'b0101010000000000000000100000000,
31'b0000000100000001100000000000000,
31'b0001100000000000100100000000000,
31'b0000000000000000000010100000001,
31'b0101010000001000000000100000000,
31'b0000000100001001100000000000000,
31'b1101000001000000000100000000000,
31'b0001000011000000011000000000000,
31'b1100000000100001000000010000000,
31'b0010000010000000110000000100000,
31'b0011000000000000010000100000000,
31'b0001000000000000000110001000000,
31'b0011000000000100010000100000000,
31'b1100000000000000000100000011000,
31'b0010100000001000000011000000000,
31'b0000000100000000001010000000010,
31'b0101010000100000000000100000000,
31'b0000001000000000011000100000000,
31'b0010100000000000000011000000000,
31'b0000000000000000110000000010000,
31'b1000001000000011000010000000000,
31'b1000001000000001000010000000000,
31'b0100011100000000000000000000000,
31'b0100011100000010000000000000000,
31'b0100011100000100000000000000000,
31'b1001000000100000100000000000001,
31'b1100000010000000000000000001100,
31'b0010000010000001000000100001000,
31'b0000001010000001000000000100000,
31'b0001000000000001001000000010000,
31'b0010001000000001000000000010000,
31'b1000100000000100000001000010000,
31'b1010000000000000110010000000000,
31'b1000100000000000000001000010000,
31'b0010001000001001000000000010000,
31'b1100110000000000000000001000000,
31'b0010001100100000010000000000000,
31'b1100000000000000101000000000100,
31'b0101000000000000100001000001000,
31'b0001000100000000011000000000000,
31'b1001000000000010100000000000001,
31'b1001000000000000100000000000001,
31'b1100010000000000100010000000000,
31'b0001000100001000011000000000000,
31'b0010100010000000000000100000100,
31'b1100100010000001000000000000000,
31'b0010001000100001000000000010000,
31'b0001000100010000011000000000000,
31'b1010000000000000000000100010001,
31'b1001000000010000100000000000001,
31'b0010000000000000000010100000010,
31'b0000010100000000000010010000000,
31'b0010001100000000010000000000000,
31'b0010010000000000000000101001000,
31'b0000000000000001001000000001000,
31'b0000010000100000100000001000000,
31'b0000010010000000000000000000110,
31'b0000100000100000001000000000100,
31'b1000010000000000000000010100000,
31'b1010000000000000000100001001000,
31'b1000010000000100000000010100000,
31'b0101100000010000000000000000001,
31'b0000110000000000000010000000000,
31'b0000110000000010000010000000000,
31'b0000110000000100000010000000000,
31'b0000000010000001100000000000000,
31'b0001000000000001000000100100000,
31'b0101100000000100000000000000001,
31'b0101100000000010000000000000001,
31'b0101100000000000000000000000001,
31'b0000010000000010100000001000000,
31'b0000010000000000100000001000000,
31'b0000100000000010001000000000100,
31'b0000100000000000001000000000100,
31'b1000010000100000000000010100000,
31'b0000010000001000100000001000000,
31'b0110100000000000010010000000000,
31'b0100000000000000100001000010000,
31'b0000110000100000000010000000000,
31'b0000010000010000100000001000000,
31'b0000110000100100000010000000000,
31'b0000100000010000001000000000100,
31'b0011101000000000000000000000100,
31'b0000010101000000000010010000000,
31'b1001001000000000000000000100001,
31'b1001000000000001000001000000100,
31'b1100000000001000000000000001100,
31'b0010000000010000000011010000000,
31'b0000010001000000000000000000110,
31'b0000000001010001100000000000000,
31'b1100000000000000000000000001100,
31'b0010000000000001000000100001000,
31'b0000001000000001000000000100000,
31'b0000000000000000000001000000101,
31'b0010001010000001000000000010000,
31'b0010000000000000000011010000000,
31'b0000011000000000010001000000000,
31'b0000000001000001100000000000000,
31'b1100000000010000000000000001100,
31'b0010000000010001000000100001000,
31'b0000001000010001000000000100000,
31'b0000000001001001100000000000000,
31'b1101000100000000000100000000000,
31'b0001000110000000011000000000000,
31'b0010100000001000000000100000100,
31'b1100100000001001000000000000000,
31'b1000000000000000000000100100001,
31'b1100100000000101000000000000000,
31'b0010100000000000000000100000100,
31'b1100100000000001000000000000000,
31'b1001000000000000001000000001001,
31'b0001000000000000100100010000000,
31'b0101000000000010001001000000000,
31'b0101000000000000001001000000000,
31'b1100000000000000001000001000010,
31'b0001010000000000001000001010000,
31'b0010100000010000000000100000100,
31'b1100100000010001000000000000000,
31'b0000010000000100000000000000110,
31'b0000000000010101100000000000000,
31'b0000010000000000000000000000110,
31'b0000000000010001100000000000000,
31'b1100000001000000000000000001100,
31'b0010000100000000100001001000000,
31'b0000010000001000000000000000110,
31'b0000000001000000000001000000101,
31'b0000110010000000000010000000000,
31'b0000000000000101100000000000000,
31'b0000000000000011100000000000000,
31'b0000000000000001100000000000000,
31'b0001100100000000100100000000000,
31'b0000000100000000000010100000001,
31'b0000010000000000000100000100001,
31'b0000000000001001100000000000000,
31'b0000100000010000100000000001100,
31'b0000010010000000100000001000000,
31'b0000100000000001000010001000000,
31'b0000100010000000001000000000100,
31'b1100000000000000010000010010000,
31'b0001010000000000010000010000010,
31'b0011001000000000000010000000010,
31'b1100100001000001000000000000000,
31'b0000100000000000100000000001100,
31'b0000000000000000001010000000010,
31'b0000010000000000001000001001000,
31'b0000000000100001100000000000000,
31'b0110000000000000010000000000110,
31'b0000000100000000110000000010000,
31'b1000000000000010001000000010001,
31'b1000000000000000001000000010001,
31'b0100100000000000000000000000000,
31'b0100100000000010000000000000000,
31'b0100100000000100000000000000000,
31'b0100100000000110000000000000000,
31'b0100100000001000000000000000000,
31'b0100100000001010000000000000000,
31'b0100100000001100000000000000000,
31'b0101000100000001000100000000000,
31'b0100100000010000000000000000000,
31'b0100100000010010000000000000000,
31'b0100100000010100000000000000000,
31'b0100100000010110000000000000000,
31'b1000000001100000100000000000000,
31'b1100001100000000000000001000000,
31'b1110000000000000000100000000010,
31'b0011010000000000000100000010000,
31'b0100100000100000000000000000000,
31'b1000001000000000000000000100000,
31'b1010000000000000000000100001000,
31'b1000001000000100000000000100000,
31'b1000000001010000100000000000000,
31'b1000001000001000000000000100000,
31'b1010000000001000000000100001000,
31'b1000001000001100000000000100000,
31'b1000000001001000100000000000000,
31'b1000001000010000000000000100000,
31'b1010000000010000000000100001000,
31'b1001000000000000100000000011000,
31'b1000000001000000100000000000000,
31'b1000000001000010100000000000000,
31'b1000000001000100100000000000000,
31'b1010001010000000000000000010000,
31'b0100100001000000000000000000000,
31'b0100100001000010000000000000000,
31'b0100100001000100000000000000000,
31'b0100100001000110000000000000000,
31'b1000000000110000100000000000000,
31'b1000100000000000000010001000000,
31'b1000110000000000000000000001010,
31'b1000100000000100000010001000000,
31'b0000001100000000000010000000000,
31'b0000000000000000000000011100000,
31'b0000000000000000010000100000010,
31'b0000000000000100000000011100000,
31'b1000000000100000100000000000000,
31'b1000000000100010100000000000000,
31'b1000000000100100100000000000000,
31'b1000000010000000000000001000110,
31'b1000000000011000100000000000000,
31'b1000001001000000000000000100000,
31'b1010000001000000000000100001000,
31'b1000001001000100000000000100000,
31'b1000000000010000100000000000000,
31'b0100000100000000000000010000000,
31'b1000000000010100100000000000000,
31'b1000000010000000001000000001000,
31'b1000000000001000100000000000000,
31'b1000000000001010100000000000000,
31'b1000000000001100100000000000000,
31'b1001000010000000000000100100000,
31'b1000000000000000100000000000000,
31'b1000000000000010100000000000000,
31'b1000000000000100100000000000000,
31'b1000000000000110100000000000000,
31'b0100100010000000000000000000000,
31'b0100100010000010000000000000000,
31'b0100100010000100000000000000000,
31'b0100100010000110000000000000000,
31'b0100100010001000000000000000000,
31'b0100100010001010000000000000000,
31'b0100100010001100000000000000000,
31'b1000001000000000010001001000000,
31'b0100100010010000000000000000000,
31'b0100100010010010000000000000000,
31'b0100000000000000000010000000110,
31'b0100100000000000101000000001000,
31'b1100000000000000000000000010101,
31'b0010000000000100011000000000010,
31'b0110100000000000000000000110000,
31'b0010000000000000011000000000010,
31'b1001000000000000001000000010000,
31'b1000001010000000000000000100000,
31'b1010000010000000000000100001000,
31'b1000001010000100000000000100000,
31'b1001000000001000001000000010000,
31'b1000001010001000000000000100000,
31'b1001001000000000100000100000000,
31'b1000000001000000001000000001000,
31'b1001000000010000001000000010000,
31'b1010000000000000101000100000000,
31'b0100110000000001000000001000000,
31'b1010001000001000000000000010000,
31'b1000000011000000100000000000000,
31'b1010001000000100000000000010000,
31'b1010001000000010000000000010000,
31'b1010001000000000000000000010000,
31'b0100100011000000000000000000000,
31'b0110010000000000000001010000000,
31'b0100100011000100000000000000000,
31'b1000000000101000001000000001000,
31'b1000100000000001001000000000100,
31'b1000100010000000000010001000000,
31'b1000010000000001100000001000000,
31'b1000000000100000001000000001000,
31'b0001000000000000000001000000100,
31'b0001000000000010000001000000100,
31'b0001000000000100000001000000100,
31'b1001000000100000000000100100000,
31'b1000000010100000100000000000000,
31'b1000000010100010100000000000000,
31'b1000000010100100100000000000000,
31'b1000000000000000000000001000110,
31'b1001000001000000001000000010000,
31'b1000001011000000000000000100000,
31'b1010000000000000100000000110000,
31'b1000000000001000001000000001000,
31'b1000000010010000100000000000000,
31'b1000000000000100001000000001000,
31'b1000000000000010001000000001000,
31'b1000000000000000001000000001000,
31'b1000000010001000100000000000000,
31'b1001000000000100000000100100000,
31'b1001000000000010000000100100000,
31'b1001000000000000000000100100000,
31'b1000000010000000100000000000000,
31'b1000000010000010100000000000000,
31'b1000000010000100100000000000000,
31'b0000000000000000010001010000000,
31'b0100100100000000000000000000000,
31'b0100100100000010000000000000000,
31'b0100100100000100000000000000000,
31'b0101000000001001000100000000000,
31'b0100100100001000000000000000000,
31'b0000000000000000100010000100000,
31'b0101000000000011000100000000000,
31'b0101000000000001000100000000000,
31'b0000001001000000000010000000000,
31'b1000100000000000100000010000000,
31'b0000100010000000010001000000000,
31'b1000100000000100100000010000000,
31'b0000100000100000000000001100000,
31'b1100001000000000000000001000000,
31'b0000100010001000010001000000000,
31'b1100001000000100000000001000000,
31'b1000000000000000000010011000000,
31'b1000001100000000000000000100000,
31'b1010000100000000000000100001000,
31'b1000010000000000000000010001010,
31'b0100000001000010000000010000000,
31'b0100000001000000000000010000000,
31'b0100100000000001010000000010000,
31'b0100000001000100000000010000000,
31'b0000100000001000000000001100000,
31'b1000100000100000100000010000000,
31'b0000100010100000010001000000000,
31'b0010010000000000000000000011100,
31'b0000100000000000000000001100000,
31'b0100000001010000000000010000000,
31'b0000100000000100000000001100000,
31'b0100000001010100000000010000000,
31'b0000001000010000000010000000000,
31'b0100000000101000000000010000000,
31'b0101000000000000010000000000100,
31'b0101000000000010010000000000100,
31'b0100000000100010000000010000000,
31'b0100000000100000000000010000000,
31'b0101000000001000010000000000100,
31'b0100000000100100000000010000000,
31'b0000001000000000000010000000000,
31'b0000001000000010000010000000000,
31'b0000001000000100000010000000000,
31'b0010010000000000010000010000000,
31'b0000001000001000000010000000000,
31'b0100000000110000000000010000000,
31'b0000001000001100000010000000000,
31'b0101011000000000000000000000001,
31'b0100000000001010000000010000000,
31'b0100000000001000000000010000000,
31'b0101000000100000010000000000100,
31'b0100000000001100000000010000000,
31'b0100000000000010000000010000000,
31'b0100000000000000000000010000000,
31'b0100000000000110000000010000000,
31'b0100000000000100000000010000000,
31'b0000001000100000000010000000000,
31'b0100000000011000000000010000000,
31'b0000001000100100000010000000000,
31'b0110000000000000000010000000101,
31'b1000000100000000100000000000000,
31'b0100000000010000000000010000000,
31'b0000000000000000011000000000001,
31'b0100000000010100000000010000000,
31'b0100100110000000000000000000000,
31'b0100100110000010000000000000000,
31'b0001000000000000000010100000000,
31'b0001000000000010000010100000000,
31'b0100100110001000000000000000000,
31'b0100010000000000000000100000001,
31'b0001000000001000000010100000000,
31'b0101000010000001000100000000000,
31'b0000100000000100010001000000000,
31'b1010001000000001010000000000000,
31'b0000100000000000010001000000000,
31'b0010000000000000100010000010000,
31'b0000100010100000000000001100000,
31'b1100001010000000000000001000000,
31'b0000100000001000010001000000000,
31'b0010000100000000011000000000010,
31'b1001000100000000001000000010000,
31'b1000001110000000000000000100000,
31'b0010100000000000000000001010000,
31'b0010100000000010000000001010000,
31'b0110110000000000000001000000000,
31'b0100000011000000000000010000000,
31'b0010100000001000000000001010000,
31'b1100011000000001000000000000000,
31'b0000100010001000000000001100000,
31'b0010000000000100010000100000001,
31'b0000100000100000010001000000000,
31'b0010000000000000010000100000001,
31'b0000100010000000000000001100000,
31'b0101010000000000000100001000000,
31'b0000100010000100000000001100000,
31'b1100000001000000000100000000001,
31'b0100000000000000000001100000010,
31'b0100000010101000000000010000000,
31'b0001000001000000000010100000000,
31'b1001000000000000001100000000100,
31'b0100000010100010000000010000000,
31'b0100000010100000000000010000000,
31'b0011000000000001000000001000100,
31'b1101000000000000000000101000000,
31'b0000001010000000000010000000000,
31'b0000001010000010000010000000000,
31'b0000100001000000010001000000000,
31'b0010010010000000010000010000000,
31'b0000001010001000000010000000000,
31'b0100001000000001000100100000000,
31'b0000101000000000000100000100001,
31'b1100000000100000000100000000001,
31'b0100000010001010000000010000000,
31'b0100000010001000000000010000000,
31'b0010100001000000000000001010000,
31'b1100000000000000000000000100110,
31'b0100000010000010000000010000000,
31'b0100000010000000000000010000000,
31'b1100000000000000110001000000000,
31'b1000000100000000001000000001000,
31'b0000001010100000000010000000000,
31'b0100000010011000000000010000000,
31'b0000101000000000001000001001000,
31'b1100000000001000000100000000001,
31'b0000000000000000000101000001000,
31'b0100000010010000000000010000000,
31'b0000000010000000011000000000001,
31'b1100000000000000000100000000001,
31'b0100101000000000000000000000000,
31'b1000000000100000000000000100000,
31'b0000000000000000000001100000100,
31'b1000000000100100000000000100000,
31'b0000000000000000100000011000000,
31'b1000000000101000000000000100000,
31'b0000000000001000000001100000100,
31'b1000000010000000010001001000000,
31'b0000000101000000000010000000000,
31'b1000000000110000000000000100000,
31'b0000000101000100000010000000000,
31'b1000010100000000000001000010000,
31'b0000000101001000000010000000000,
31'b1100000100000000000000001000000,
31'b0000000101001100000010000000000,
31'b1100000100000100000000001000000,
31'b1000000000000010000000000100000,
31'b1000000000000000000000000100000,
31'b1000000000000110000000000100000,
31'b1000000000000100000000000100000,
31'b1000000000001010000000000100000,
31'b1000000000001000000000000100000,
31'b1001000010000000100000100000000,
31'b1000000000001100000000000100000,
31'b1000000000010010000000000100000,
31'b1000000000010000000000000100000,
31'b1000000001000000001000100010000,
31'b1000000000010100000000000100000,
31'b1000001001000000100000000000000,
31'b0000100000000000000010010000000,
31'b1010000010000010000000000010000,
31'b1010000010000000000000000010000,
31'b0000000100010000000010000000000,
31'b1000000001100000000000000100000,
31'b0000000100010100000010000000000,
31'b1000000001100100000000000100000,
31'b0000000100011000000010000000000,
31'b1000101000000000000010001000000,
31'b0010000100000000000000010000101,
31'b0011000000000001000000000010001,
31'b0000000100000000000010000000000,
31'b0000000100000010000010000000000,
31'b0000000100000100000010000000000,
31'b0000010000000000000100100100000,
31'b0000000100001000000010000000000,
31'b0100100000000000100000000100000,
31'b0000000100001100000010000000000,
31'b0101010100000000000000000000001,
31'b1000000001000010000000000100000,
31'b1000000001000000000000000100000,
31'b1000000001000110000000000100000,
31'b1000000001000100000000000100000,
31'b1000001000010000100000000000000,
31'b1000000001001000000000000100000,
31'b1001000000000000000000000111000,
31'b1000001010000000001000000001000,
31'b0000000100100000000010000000000,
31'b1000000001010000000000000100000,
31'b1000000000000000001000100010000,
31'b1000000001010100000000000100000,
31'b1000001000000000100000000000000,
31'b1000001000000010100000000000000,
31'b1000001000000100100000000000000,
31'b1010000011000000000000000010000,
31'b0001000000000000010000000000010,
31'b1000000010100000000000000100000,
31'b0001000000000100010000000000010,
31'b1000000010100100000000000100000,
31'b0001000000001000010000000000010,
31'b1000000010101000000000000100000,
31'b1001000000100000100000100000000,
31'b1000000000000000010001001000000,
31'b0001000000010000010000000000010,
31'b1010000100000001010000000000000,
31'b0101100001000000000000100000000,
31'b1010000000101000000000000010000,
31'b0001010001000000100100000000000,
31'b1100000110000000000000001000000,
31'b1010000000100010000000000010000,
31'b1010000000100000000000000010000,
31'b1000000010000010000000000100000,
31'b1000000010000000000000000100000,
31'b1001000000001000100000100000000,
31'b1000000010000100000000000100000,
31'b1001000000000100100000100000000,
31'b1000000010001000000000000100000,
31'b1001000000000000100000100000000,
31'b0000000000000000000000010000110,
31'b1011000001000000000000000001000,
31'b1000000010010000000000000100000,
31'b1010000000001010000000000010000,
31'b1010000000001000000000000010000,
31'b1010000000000110000000000010000,
31'b1010000000000100000000000010000,
31'b1010000000000010000000000010000,
31'b1010000000000000000000000010000,
31'b0001000001000000010000000000010,
31'b1000000011100000000000000100000,
31'b0100000000000000010011000000000,
31'b0110100000000000100000000010000,
31'b0001010000010000100100000000000,
31'b0010010000000000000100100010000,
31'b0100100000000000001000000101000,
31'b0010000000000000001001000000100,
31'b0000000110000000000010000000000,
31'b0001000000000001000000000100001,
31'b0101100000000000000000100000000,
31'b0101100000000010000000100000000,
31'b0001010000000000100100000000000,
31'b0100100010000000100000000100000,
31'b0101100000001000000000100000000,
31'b1010000001100000000000000010000,
31'b1011000000010000000000000001000,
31'b1000000011000000000000000100000,
31'b0100100000000000000100001000001,
31'b1000001000001000001000000001000,
31'b1010000000000000001000100100000,
31'b1000001000000100001000000001000,
31'b1001000001000000100000100000000,
31'b1000001000000000001000000001000,
31'b1011000000000000000000000001000,
31'b1011000000000010000000000001000,
31'b1011000000000100000000000001000,
31'b1010000001001000000000000010000,
31'b1000001010000000100000000000000,
31'b1010000001000100000000000010000,
31'b1010000001000010000000000010000,
31'b1010000001000000000000000010000,
31'b0000000001010000000010000000000,
31'b1000000100100000000000000100000,
31'b0000000100000000000001100000100,
31'b1000010000010000000001000010000,
31'b0000000100000000100000011000000,
31'b1100000000010000000000001000000,
31'b0010000001000000000000010000101,
31'b1100000000010100000000001000000,
31'b0000000001000000000010000000000,
31'b0000000001000010000010000000000,
31'b0000000001000100000010000000000,
31'b1000010000000000000001000010000,
31'b0000000001001000000010000000000,
31'b1100000000000000000000001000000,
31'b0000000001001100000010000000000,
31'b1100000000000100000000001000000,
31'b1000000100000010000000000100000,
31'b1000000100000000000000000100000,
31'b1000010000000000000110100000000,
31'b1000000100000100000000000100000,
31'b1100100000000000100010000000000,
31'b1000000100001000000000000100000,
31'b0010010010000000000000100000100,
31'b1100010010000001000000000000000,
31'b0000000001100000000010000000000,
31'b1000000100010000000000000100000,
31'b0000000001100100000010000000000,
31'b1000010000100000000001000010000,
31'b0000101000000000000000001100000,
31'b1100000000100000000000001000000,
31'b0000101000000100000000001100000,
31'b1100000000100100000000001000000,
31'b0000000000010000000010000000000,
31'b0000000000010010000010000000000,
31'b0000000000010100000010000000000,
31'b0000010000100000001000000000100,
31'b0000000000011000000010000000000,
31'b0100001000100000000000010000000,
31'b0010000000000000000000010000101,
31'b0101010000010000000000000000001,
31'b0000000000000000000010000000000,
31'b0000000000000010000010000000000,
31'b0000000000000100000010000000000,
31'b0000000000000110000010000000000,
31'b0000000000001000000010000000000,
31'b0000000000001010000010000000000,
31'b0000000000001100000010000000000,
31'b0101010000000000000000000000001,
31'b0000000000110000000010000000000,
31'b0000100000000000100000001000000,
31'b0000010000000010001000000000100,
31'b0000010000000000001000000000100,
31'b0100001000000010000000010000000,
31'b0100001000000000000000010000000,
31'b0110010000000000010010000000000,
31'b0100001000000100000000010000000,
31'b0000000000100000000010000000000,
31'b0000000000100010000010000000000,
31'b0000000000100100000010000000000,
31'b0000010000010000001000000000100,
31'b0000000000101000000010000000000,
31'b0100001000010000000000010000000,
31'b0000001000000000011000000000001,
31'b0101010000100000000000000000001,
31'b0001000100000000010000000000010,
31'b1010000000010001010000000000000,
31'b0001001000000000000010100000000,
31'b0001001000000010000010100000000,
31'b0001000100001000010000000000010,
31'b1100000010010000000000001000000,
31'b0010010000100000000000100000100,
31'b1100010000100001000000000000000,
31'b0000000011000000000010000000000,
31'b1010000000000001010000000000000,
31'b0000101000000000010001000000000,
31'b1010000000000101010000000000000,
31'b0000000011001000000010000000000,
31'b1100000010000000000000001000000,
31'b0000101000001000010001000000000,
31'b1100000010000100000000001000000,
31'b1001000000000001000010000000001,
31'b1000000110000000000000000100000,
31'b0010101000000000000000001010000,
31'b1100010000001001000000000000000,
31'b0010010000000100000000100000100,
31'b1100010000000101000000000000000,
31'b0010010000000000000000100000100,
31'b1100010000000001000000000000000,
31'b0000000011100000000010000000000,
31'b1010000000100001010000000000000,
31'b0000101000100000010001000000000,
31'b1100000000000000010001000100000,
31'b0000101010000000000000001100000,
31'b1100000010100000000000001000000,
31'b1100000000000000100000000000110,
31'b1010000100000000000000000010000,
31'b0000000010010000000010000000000,
31'b0000000010010010000010000000000,
31'b0000100000000000000000000000110,
31'b0000100000000010000000000000110,
31'b0000000010011000000010000000000,
31'b0100001010100000000000010000000,
31'b0010000000000000000010000110000,
31'b0010000100000000001001000000100,
31'b0000000010000000000010000000000,
31'b0000000010000010000010000000000,
31'b0000000010000100000010000000000,
31'b0000110000000001100000000000000,
31'b0000000010001000000010000000000,
31'b0100000000000001000100100000000,
31'b0000100000000000000100000100001,
31'b0101010010000000000000000000001,
31'b0000000010110000000010000000000,
31'b0000000000000001000000000001010,
31'b0000100000100000000000000000110,
31'b0000010010000000001000000000100,
31'b0100001010000010000000010000000,
31'b0100001010000000000000010000000,
31'b0010010001000000000000100000100,
31'b1100010001000001000000000000000,
31'b0000000010100000000010000000000,
31'b0000000010100010000010000000000,
31'b0000100000000000001000001001000,
31'b0000110000100001100000000000000,
31'b0000001000000000000101000001000,
31'b0100001010010000000000010000000,
31'b0000100000100000000100000100001,
31'b1100001000000000000100000000001,
31'b0100110000000000000000000000000,
31'b0100110000000010000000000000000,
31'b0100110000000100000000000000000,
31'b0100110000000110000000000000000,
31'b0100110000001000000000000000000,
31'b0100110000001010000000000000000,
31'b0000000000000000100100100000000,
31'b0001100000000000000010000000001,
31'b0100110000010000000000000000000,
31'b0100110000010010000000000000000,
31'b0100110000010100000000000000000,
31'b1001000000000000000000010100001,
31'b1100000000000000010000100001000,
31'b0011000000000100000100000010000,
31'b0010100000100000010000000000000,
31'b0011000000000000000100000010000,
31'b1000000000000000010100000000010,
31'b1000011000000000000000000100000,
31'b1010010000000000000000100001000,
31'b1000011000000100000000000100000,
31'b1000010001010000100000000000000,
31'b1000011000001000000000000100000,
31'b0010100000010000010000000000000,
31'b0010100000010010010000000000000,
31'b1000010001001000100000000000000,
31'b1000011000010000000000000100000,
31'b0100000000000000100000000001010,
31'b0100100000000000001010000000100,
31'b1000010001000000100000000000000,
31'b1000010001000010100000000000000,
31'b0010100000000000010000000000000,
31'b0010100000000010010000000000000,
31'b0100110001000000000000000000000,
31'b0110000010000000000001010000000,
31'b1110000000000000110000000000000,
31'b0010000100010000010000010000000,
31'b1000100000000100000000000001010,
31'b1000110000000000000010001000000,
31'b1000100000000000000000000001010,
31'b1000100000000010000000000001010,
31'b0010000000000000000100000001000,
31'b0010000000000010000100000001000,
31'b0010000000000100000100000001000,
31'b0010000100000000010000010000000,
31'b1000010000100000100000000000000,
31'b1000010000100010100000000000000,
31'b1000100000010000000000000001010,
31'b0101001100000000000000000000001,
31'b1000010000011000100000000000000,
31'b1000011001000000000000000100000,
31'b0001000100000000000010010000001,
31'b0000001100000000001000000000100,
31'b1000010000010000100000000000000,
31'b1000000000000001000000000000110,
31'b1000100000100000000000000001010,
31'b1000010010000000001000000001000,
31'b1000010000001000100000000000000,
31'b1000010000001010100000000000000,
31'b1100100000000000000100100000000,
31'b0010100000000001000100000000100,
31'b1000010000000000100000000000000,
31'b1000010000000010100000000000000,
31'b1000010000000100100000000000000,
31'b1000100010000001000010000000000,
31'b0100110010000000000000000000000,
31'b0001000000000000000100000100000,
31'b0100110010000100000000000000000,
31'b0100000000000001100010000000000,
31'b0100110010001000000000000000000,
31'b0100000100000000000000100000001,
31'b0000100100000001000000000100000,
31'b0100000100000100000000100000001,
31'b0100110010010000000000000000000,
31'b0100000000000000000000001001100,
31'b1000000100000001000010010000000,
31'b1001000000000000000010000010100,
31'b1000000001000000000010000001100,
31'b0001000000000000000000000000111,
31'b0010100010100000010000000000000,
31'b0011000010000000000100000010000,
31'b0100000000000010001000000000010,
31'b0100000000000000001000000000010,
31'b0100100000010001000000001000000,
31'b0100000000000100001000000000010,
31'b0110100100000000000001000000000,
31'b0100000000001000001000000000010,
31'b0010100010010000010000000000000,
31'b1100001100000001000000000000000,
31'b0100100000000101000000001000000,
31'b0100000000010000001000000000010,
31'b0100100000000001000000001000000,
31'b0100100000000011000000001000000,
31'b1000010011000000100000000000000,
31'b0101000100000000000100001000000,
31'b0010100010000000010000000000000,
31'b1010011000000000000000000010000,
31'b0110000000000010000001010000000,
31'b0110000000000000000001010000000,
31'b1010000000000000000000010001001,
31'b0010000000000000101100000000000,
31'b1000000000010000000010000001100,
31'b0110000000001000000001010000000,
31'b1000000000000001100000001000000,
31'b1000010000100000001000000001000,
31'b0010000010000000000100000001000,
31'b0110000000010000000001010000000,
31'b0010000010000100000100000001000,
31'b0010000110000000010000010000000,
31'b1000000000000000000010000001100,
31'b1000100000000000101000000000010,
31'b1000000000010001100000001000000,
31'b1000100000100001000010000000000,
31'b0100100000000000000000110000001,
31'b0100000001000000001000000000010,
31'b0000000000000011000000010100000,
31'b0000000000000001000000010100000,
31'b1000010010010000100000000000000,
31'b1000010000000100001000000001000,
31'b1000010000000010001000000001000,
31'b1000010000000000001000000001000,
31'b1001000100000000000110000000000,
31'b0100000001010000001000000000010,
31'b0100100001000001000000001000000,
31'b0000100000000000011000100000000,
31'b1000010010000000100000000000000,
31'b1000100000000101000010000000000,
31'b1000100000000011000010000000000,
31'b1000100000000001000010000000000,
31'b0100110100000000000000000000000,
31'b0100110100000010000000000000000,
31'b0101000000000000100000000100001,
31'b1000001000010000000001000010000,
31'b0100110100001000000000000000000,
31'b0100000010000000000000100000001,
31'b0000100010000001000000000100000,
31'b0101010000000001000100000000000,
31'b0010100000000001000000000010000,
31'b1000110000000000100000010000000,
31'b1000001000000010000001000010000,
31'b1000001000000000000001000010000,
31'b0011000001100000000000000000100,
31'b1100011000000000000000001000000,
31'b0010100100100000010000000000000,
31'b1100000000000000000100110000000,
31'b1000010000000000000010011000000,
31'b1000011100000000000000000100000,
31'b1000001000000000000110100000000,
31'b1000000000000000000000010001010,
31'b0110100010000000000001000000000,
31'b0100010001000000000000010000000,
31'b0010100100010000010000000000000,
31'b1100001010000001000000000000000,
31'b0011000001001000000000000000100,
31'b0011000000000001010100000000000,
31'b0100100000000000000001000110000,
31'b0010000000000000000000000011100,
31'b0011000001000000000000000000100,
31'b0101000010000000000100001000000,
31'b0010100100000000010000000000000,
31'b0010100100000010010000000000000,
31'b0110000000000000001000000000001,
31'b0110000000000010001000000000001,
31'b0110000000000100001000000000001,
31'b0010000000010000010000010000000,
31'b0110000000001000001000000000001,
31'b0100010000100000000000010000000,
31'b1000100100000000000000000001010,
31'b0101001000010000000000000000001,
31'b0000011000000000000010000000000,
31'b0010000000000100010000010000000,
31'b0010000000000010010000010000000,
31'b0010000000000000010000010000000,
31'b0011000000100000000000000000100,
31'b0101001000000100000000000000001,
31'b0101001000000010000000000000001,
31'b0101001000000000000000000000001,
31'b0110000000100000001000000000001,
31'b0100010000001000000000010000000,
31'b0001000000000000000010010000001,
31'b0000001000000000001000000000100,
31'b0100010000000010000000010000000,
31'b0100010000000000000000010000000,
31'b0110001000000000010010000000000,
31'b0100010000000100000000010000000,
31'b0011000000001000000000000000100,
31'b0101000000000000011010000000000,
31'b0011000000001100000000000000100,
31'b0010000000100000010000010000000,
31'b0011000000000000000000000000100,
31'b0100010000010000000000010000000,
31'b0011000000000100000000000000100,
31'b0101001000100000000000000000001,
31'b0100110110000000000000000000000,
31'b0100000000001000000000100000001,
31'b0001010000000000000010100000000,
31'b0100000100000001100010000000000,
31'b0100000000000010000000100000001,
31'b0100000000000000000000100000001,
31'b0000100000000001000000000100000,
31'b0100000000000100000000100000001,
31'b1010000001000000100001000000000,
31'b0100000100000000000000001001100,
31'b1000000000000001000010010000000,
31'b1000001010000000000001000010000,
31'b0100100000000000010000001010000,
31'b0100000000010000000000100000001,
31'b0000100000010001000000000100000,
31'b0100000001000001000000011000000,
31'b0110100000001000000001000000000,
31'b0100000100000000001000000000010,
31'b0010110000000000000000001010000,
31'b1100001000001001000000000000000,
31'b0110100000000000000001000000000,
31'b0000000000000000000000000101100,
31'b0010001000000000000000100000100,
31'b1100001000000001000000000000000,
31'b1001000001000000000110000000000,
31'b0001000000000000001000100000100,
31'b1100000000000000000101000000010,
31'b0010010000000000010000100000001,
31'b0110100000010000000001000000000,
31'b0101000000000000000100001000000,
31'b0010100110000000010000000000000,
31'b1100001000010001000000000000000,
31'b1010000000010000100001000000000,
31'b1010000000000000010100000000001,
31'b0001010001000000000010100000000,
31'b0010000100000000101100000000000,
31'b0100100000000000001000010000010,
31'b0100000001000000000000100000001,
31'b0000100001000001000000000100000,
31'b0100000001000100000000100000001,
31'b1010000000000000100001000000000,
31'b1010000000000010100001000000000,
31'b1010000000000100100001000000000,
31'b0010000010000000010000010000000,
31'b1010000000001000100001000000000,
31'b0100000001010000000000100000001,
31'b0100000000000011000000011000000,
31'b0100000000000001000000011000000,
31'b1001000000010000000110000000000,
31'b0100010010001000000000010000000,
31'b0001000000000000000000000110100,
31'b0000001010000000001000000000100,
31'b0110100001000000000001000000000,
31'b0100010010000000000000010000000,
31'b0011100000000000000010000000010,
31'b1100001001000001000000000000000,
31'b1001000000000000000110000000000,
31'b1001000000000010000110000000000,
31'b1100000000000001100000000100000,
31'b0010000010100000010000010000000,
31'b0011000010000000000000000000100,
31'b0101000001000000000100001000000,
31'b0011000010000100000000000000100,
31'b1100010000000000000100000000001,
31'b0000000000000000001100000010000,
31'b1000010000100000000000000100000,
31'b0000010000000000000001100000100,
31'b1000010000100100000000000100000,
31'b0000010000000000100000011000000,
31'b1010000000000001000000001010000,
31'b0000100000000000001000010000100,
31'b0001101000000000000010000000001,
31'b0000010101000000000010000000000,
31'b1000010000110000000000000100000,
31'b1000000100000010000001000010000,
31'b1000000100000000000001000010000,
31'b0001000100000000000000001010010,
31'b1100010100000000000000001000000,
31'b0010101000100000010000000000000,
31'b1110000000000000010000000100000,
31'b1000010000000010000000000100000,
31'b1000010000000000000000000100000,
31'b1000010000000110000000000100000,
31'b1000010000000100000000000100000,
31'b1000010000001010000000000100000,
31'b1000010000001000000000000100000,
31'b0010101000010000010000000000000,
31'b1100000110000001000000000000000,
31'b1000010000010010000000000100000,
31'b1000010000010000000000000100000,
31'b0101100000000000000000010000001,
31'b1000010000010100000000000100000,
31'b1000011001000000100000000000000,
31'b1000000000000001010001000000000,
31'b0010101000000000010000000000000,
31'b1010010010000000000000000010000,
31'b0000010100010000000010000000000,
31'b1000010001100000000000000100000,
31'b0000010100010100000010000000000,
31'b0000000100100000001000000000100,
31'b0001000100000000011000010000000,
31'b0010000010000000000100100010000,
31'b1001000000000000100000010000001,
31'b0001000000000000001100000001000,
31'b0000010100000000000010000000000,
31'b0000010100000010000010000000000,
31'b0000010100000100000010000000000,
31'b0000000000000000000100100100000,
31'b0001000010000000100100000000000,
31'b0101000100000100000000000000001,
31'b0101000100000010000000000000001,
31'b0101000100000000000000000000001,
31'b1000010001000010000000000100000,
31'b1000010001000000000000000100000,
31'b0000000100000010001000000000100,
31'b0000000100000000001000000000100,
31'b1000011000010000100000000000000,
31'b1000010001001000000000000100000,
31'b0110000100000000010010000000000,
31'b0100000000000000000000000101010,
31'b1000000000000000000101000000100,
31'b1000010001010000000000000100000,
31'b1000010000000000001000100010000,
31'b0000000100010000001000000000100,
31'b1000011000000000100000000000000,
31'b1000011000000010100000000000000,
31'b1000100000000000000001010010000,
31'b0101000100100000000000000000001,
31'b0001010000000000010000000000010,
31'b1100000000000000010000000010000,
31'b0011000000000000000100100001000,
31'b1100000000000100010000000010000,
31'b0001010000001000010000000000010,
31'b1100000000001000010000000010000,
31'b0010000100100000000000100000100,
31'b1100000100100001000000000000000,
31'b0001010000010000010000000000010,
31'b1100000000010000010000000010000,
31'b1000000000000011000000001100000,
31'b1000000000000001000000001100000,
31'b0001000001000000100100000000000,
31'b0001001000000000000000000000111,
31'b0010000000000000001100000100000,
31'b1010010000100000000000000010000,
31'b1101100000000000000100000000000,
31'b1000010010000000000000000100000,
31'b0010000100001000000000100000100,
31'b1100000100001001000000000000000,
31'b0010000100000100000000100000100,
31'b1100000100000101000000000000000,
31'b0010000100000000000000100000100,
31'b1100000100000001000000000000000,
31'b0010000001001000000011000000000,
31'b1110000000000000000001001000000,
31'b0010000000000000000000001001001,
31'b1010010000001000000000000010000,
31'b0010000001000000000011000000000,
31'b1010010000000100000000000010000,
31'b0000000000000001100000010000000,
31'b1010010000000000000000000010000,
31'b0001010001000000010000000000010,
31'b1100000001000000010000000010000,
31'b1100100000000001000000010000000,
31'b0010100000000000000000110000100,
31'b0001000000010000100100000000000,
31'b0010000000000000000100100010000,
31'b1101000000000000010000000001000,
31'b0010010000000000001001000000100,
31'b0001000000001000100100000000000,
31'b0001010000000001000000000100001,
31'b0101110000000000000000100000000,
31'b0000100100000001100000000000000,
31'b0001000000000000100100000000000,
31'b0001000000000010100100000000000,
31'b0100000000000001000010000100000,
31'b0101000110000000000000000000001,
31'b0010000000011000000011000000000,
31'b1100000000000000000000010001100,
31'b0000000100000001000010001000000,
31'b0000001000000001000000010100000,
31'b0010000000010000000011000000000,
31'b0010000000100000000100100010000,
31'b0010000101000000000000100000100,
31'b1100000101000001000000000000000,
31'b0010000000001000000011000000000,
31'b0110000000000000000000000011010,
31'b0010000001000000000000001001001,
31'b0000101000000000011000100000000,
31'b0010000000000000000011000000000,
31'b0010000000000010000011000000000,
31'b0010000000000100000011000000000,
31'b1010010001000000000000000010000,
31'b0000010001010000000010000000000,
31'b1000010100100000000000000100000,
31'b1000000000100000000110100000000,
31'b1000000000010000000001000010000,
31'b0001000001000000011000010000000,
31'b1100010000010000000000001000000,
31'b0010000010100000000000100000100,
31'b1100000010100001000000000000000,
31'b0000010001000000000010000000000,
31'b1000000000000100000001000010000,
31'b1000000000000010000001000010000,
31'b1000000000000000000001000010000,
31'b0001000000000000000000001010010,
31'b1100010000000000000000001000000,
31'b1100000000000000000010000001010,
31'b1000000000001000000001000010000,
31'b1000010100000010000000000100000,
31'b1000010100000000000000000100000,
31'b1000000000000000000110100000000,
31'b0000000001000000001000000000100,
31'b0011000000000000010001000000010,
31'b1100000010000101000000000000000,
31'b0010000010000000000000100000100,
31'b1100000010000001000000000000000,
31'b0000010001100000000010000000000,
31'b1000010100010000000000000100000,
31'b1000000000100010000001000010000,
31'b1000000000100000000001000010000,
31'b0011001001000000000000000000100,
31'b1100010000100000000000001000000,
31'b0010101100000000010000000000000,
31'b1100000010010001000000000000000,
31'b0000010000010000000010000000000,
31'b0000010000010010000010000000000,
31'b0000010000010100000010000000000,
31'b0000000000100000001000000000100,
31'b0001000000000000011000010000000,
31'b0101000000010100000000000000001,
31'b0110000000100000010010000000000,
31'b0101000000010000000000000000001,
31'b0000010000000000000010000000000,
31'b0000010000000010000010000000000,
31'b0000010000000100000010000000000,
31'b0000000000000000000000001001010,
31'b0000010000001000000010000000000,
31'b0101000000000100000000000000001,
31'b0101000000000010000000000000001,
31'b0101000000000000000000000000001,
31'b0000010000110000000010000000000,
31'b0000000000000100001000000000100,
31'b0000000000000010001000000000100,
31'b0000000000000000001000000000100,
31'b0110000000000100010010000000000,
31'b0100011000000000000000010000000,
31'b0110000000000000010010000000000,
31'b0000000000001000001000000000100,
31'b0000010000100000000010000000000,
31'b0000010000100010000010000000000,
31'b0000010000100100000010000000000,
31'b0000000000010000001000000000100,
31'b0011001000000000000000000000100,
31'b0101000000100100000000000000001,
31'b0110000000010000010010000000000,
31'b0101000000100000000000000000001,
31'b0001010100000000010000000000010,
31'b1100000100000000010000000010000,
31'b0011000000000000000000001100010,
31'b1100000000101001000000000000000,
31'b1100100000000000000000000001100,
31'b1010000000000000000001000100000,
31'b0010000000100000000000100000100,
31'b1100000000100001000000000000000,
31'b0000010011000000000010000000000,
31'b1010010000000001010000000000000,
31'b1000001000000001000010010000000,
31'b1000000010000000000001000010000,
31'b0001000101000000100100000000000,
31'b1100010010000000000000001000000,
31'b0010000100000000001100000100000,
31'b1100000000110001000000000000000,
31'b0010000000001100000000100000100,
31'b1100000000001101000000000000000,
31'b0010000000001000000000100000100,
31'b1100000000001001000000000000000,
31'b0010000000000100000000100000100,
31'b1100000000000101000000000000000,
31'b0010000000000000000000100000100,
31'b1100000000000001000000000000000,
31'b0000000001000000100000000001100,
31'b0001100000000000100100010000000,
31'b0010000100000000000000001001001,
31'b1100000000011001000000000000000,
31'b0010000101000000000011000000000,
31'b1100000000010101000000000000000,
31'b0010000000010000000000100000100,
31'b1100000000010001000000000000000,
31'b0000010010010000000010000000000,
31'b0000100000010101100000000000000,
31'b0000110000000000000000000000110,
31'b0000100000010001100000000000000,
31'b0001000100010000100100000000000,
31'b1101000000000000000100010000000,
31'b0010010000000000000010000110000,
31'b1100000001100001000000000000000,
31'b0000010010000000000010000000000,
31'b0000100000000101100000000000000,
31'b0000100000000011100000000000000,
31'b0000100000000001100000000000000,
31'b0001000100000000100100000000000,
31'b0101000010000100000000000000001,
31'b0101000010000010000000000000001,
31'b0101000010000000000000000000001,
31'b0000000000010000100000000001100,
31'b0000010000000001000000000001010,
31'b0000000000000001000010001000000,
31'b0000000010000000001000000000100,
31'b0010000100010000000011000000000,
31'b1100000001000101000000000000000,
31'b0010000001000000000000100000100,
31'b1100000001000001000000000000000,
31'b0000000000000000100000000001100,
31'b0000100000000000001010000000010,
31'b0000000000010001000010001000000,
31'b0000100000100001100000000000000,
31'b0010000100000000000011000000000,
31'b0010000100000010000011000000000,
31'b0010000100000100000011000000000,
31'b1100000001010001000000000000000,
31'b0101000000000000000000000000000,
31'b0101000000000010000000000000000,
31'b0101000000000100000000000000000,
31'b0101000000000110000000000000000,
31'b0101000000001000000000000000000,
31'b0101000000001010000000000000000,
31'b0101000000001100000000000000000,
31'b0000010000000000000010000000001,
31'b0101000000010000000000000000000,
31'b0101000000010010000000000000000,
31'b0101000000010100000000000000000,
31'b0110001000001000001000000000000,
31'b0101000000011000000000000000000,
31'b0110001000000100001000000000000,
31'b0110001000000010001000000000000,
31'b0110001000000000001000000000000,
31'b0101000000100000000000000000000,
31'b0101000000100010000000000000000,
31'b0101000000100100000000000000000,
31'b0101000000100110000000000000000,
31'b0101000000101000000000000000000,
31'b0101000000101010000000000000000,
31'b0101000000101100000000000000000,
31'b0100000000000000010000010000100,
31'b0101000000110000000000000000000,
31'b0110000000000000010010000000001,
31'b0101000000110100000000000000000,
31'b1000100000000000100000000011000,
31'b0000000000000000001000000000101,
31'b0001001000000000000010010000000,
31'b0011010000000000010000000000000,
31'b0110001000100000001000000000000,
31'b0101000001000000000000000000000,
31'b0101000001000010000000000000000,
31'b0000000000000000000011000000010,
31'b0100000000001000000000000011000,
31'b1000000000000000000001000010001,
31'b1001000000000000000010001000000,
31'b0100000000000010000000000011000,
31'b0100000000000000000000000011000,
31'b0101000001010000000000000000000,
31'b0110000010000000000000000101000,
31'b0100001010000000000000100000000,
31'b0100001010000010000000100000000,
31'b1001100000100000100000000000000,
31'b1001000000010000000010001000000,
31'b0100001010001000000000100000000,
31'b0100000000010000000000000011000,
31'b0101000001100000000000000000000,
31'b0101000001100010000000000000000,
31'b0100000000000001000100010000000,
31'b0100000000101000000000000011000,
31'b1001100000010000100000000000000,
31'b1010100000000000000000100010000,
31'b0100000000100010000000000011000,
31'b0100000000100000000000000011000,
31'b1100000010000001000000000000001,
31'b0010010000000000010000000011000,
31'b0100001010100000000000100000000,
31'b0000000010000001000001000001000,
31'b1001100000000000100000000000000,
31'b1001100000000010100000000000000,
31'b1001100000000100100000000000000,
31'b0100001000000000000001010000010,
31'b0101000010000000000000000000000,
31'b0101000010000010000000000000000,
31'b0101000010000100000000000000000,
31'b0101000010000110000000000000000,
31'b0101000010001000000000000000000,
31'b0101000010001010000000000000000,
31'b0101000010001100000000000000000,
31'b0100000000000000100000100100000,
31'b0101000010010000000000000000000,
31'b0110000001000000000000000101000,
31'b0100001001000000000000100000000,
31'b0101000000000000101000000001000,
31'b0101000010011000000000000000000,
31'b1000010000000000000110010000000,
31'b1010001000000000010100000000000,
31'b1010010000000000000000000100010,
31'b1000100000000000001000000010000,
31'b1100000000000000010000000100010,
31'b1100000000000000000000111000000,
31'b0010000100000000000011000000001,
31'b1100000000000000100001000000100,
31'b0010000101000000000000001001000,
31'b1000101000000000100000100000000,
31'b0000000001000000000010110000000,
31'b1100000001000001000000000000001,
31'b0010000001000000000000100000101,
31'b0101010000000001000000001000000,
31'b0000000100000000100000101000000,
31'b0001000000000001000001000010000,
31'b0000000100000000000001010000100,
31'b0011010010000000010000000000000,
31'b0000000100001000100000101000000,
31'b0101000011000000000000000000000,
31'b0110000000010000000000000101000,
31'b0100001000010000000000100000000,
31'b0100001000010010000000100000000,
31'b1001000000000001001000000000100,
31'b1001000010000000000010001000000,
31'b0100001000011000000000100000000,
31'b0100000010000000000000000011000,
31'b0000100000000000000001000000100,
31'b0110000000000000000000000101000,
31'b0100001000000000000000100000000,
31'b0100001000000010000000100000000,
31'b0100000000000000101000000010000,
31'b0110000000001000000000000101000,
31'b0100001000001000000000100000000,
31'b0100001000001010000000100000000,
31'b1100000000010001000000000000001,
31'b0010000100001000000000001001000,
31'b0100001000110000000000100000000,
31'b0000000000010001000001000001000,
31'b0010011000000000010000100000000,
31'b0010000100000000000000001001000,
31'b0000001000000000000100000001010,
31'b0000000000000000000010110000000,
31'b1100000000000001000000000000001,
31'b0010000000000000000000100000101,
31'b0100001000100000000000100000000,
31'b0000000000000001000001000001000,
31'b1100000000001001000000000000001,
31'b0010000100010000000000001001000,
31'b0100001000101000000000100000000,
31'b0000000000010000000010110000000,
31'b0101000100000000000000000000000,
31'b0101000100000010000000000000000,
31'b0101000100000100000000000000000,
31'b0101000100000110000000000000000,
31'b0101000100001000000000000000000,
31'b0101000100001010000000000000000,
31'b0101000100001100000000000000000,
31'b0100100000000001000100000000000,
31'b0000000000000000000000100000110,
31'b1001000000000000100000010000000,
31'b0001000010000000010001000000000,
31'b1001000000000100100000010000000,
31'b0001000000100000000000001100000,
31'b1001000000001000100000010000000,
31'b1000000010000000000000110100000,
31'b0110001100000000001000000000000,
31'b0101000100100000000000000000000,
31'b0101000100100010000000000000000,
31'b0101000100100100000000000000000,
31'b1000011000000000100000000000001,
31'b0100000000000000000100000001100,
31'b0101100001000000000000010000000,
31'b1000001000000001000100000100000,
31'b1000010000000001010000000000010,
31'b0001000000001000000000001100000,
31'b1001000000100000100000010000000,
31'b1000000000001000110000000000100,
31'b1000000000000000000001000100010,
31'b0001000000000000000000001100000,
31'b0001000000000010000000001100000,
31'b1000000000000000110000000000100,
31'b1000000000001000000001000100010,
31'b0101000101000000000000000000000,
31'b0101000101000010000000000000000,
31'b0100100000000000010000000000100,
31'b0100100000000010010000000000100,
31'b1001001000000000000000010100000,
31'b1001000100000000000010001000000,
31'b0100100000001000010000000000100,
31'b0100000100000000000000000011000,
31'b0001101000000000000010000000000,
31'b1001000001000000100000010000000,
31'b0100100000010000010000000000100,
31'b1010000000000000001000010100000,
31'b0010110000100000000000000000100,
31'b0010010000000101000000000001000,
31'b1000010000100000000000000100001,
31'b0010010000000001000000000001000,
31'b0101000101100000000000000000000,
31'b0100000000000001010000000001000,
31'b1000010000000000000100000000110,
31'b1000001000000000010000000100100,
31'b0101100000000010000000010000000,
31'b0101100000000000000000010000000,
31'b1000010000010000000000000100001,
31'b0101100000000100000000010000000,
31'b0010110000001000000000000000100,
31'b1101000000000000000010000100000,
31'b1000010000001000000000000100001,
31'b1000000000000001100100000000000,
31'b0010110000000000000000000000100,
31'b0101100000010000000000010000000,
31'b1000010000000000000000000100001,
31'b1000010000000010000000000100001,
31'b0101000110000000000000000000000,
31'b0101000110000010000000000000000,
31'b0000100000000000000010100000000,
31'b0001000000000000100100000000001,
31'b0101000110001000000000000000000,
31'b1000000001000000001000010010000,
31'b0001010000000001000000000100000,
31'b0100100010000001000100000000000,
31'b0001000000000100010001000000000,
31'b1001000010000000100000010000000,
31'b0001000000000000010001000000000,
31'b0001000000000010010001000000000,
31'b1000000000000100000000110100000,
31'b1000000000000000010000001000010,
31'b1000000000000000000000110100000,
31'b1000000000000100010000001000010,
31'b1110000000000000000010000001000,
31'b0010000001001000000000001001000,
31'b0011000000000000000000001010000,
31'b0010000000000000000011000000001,
31'b0111010000000000000001000000000,
31'b0010000001000000000000001001000,
31'b0011000000001000000000001010000,
31'b0010000001000100000000001001000,
31'b0001000010001000000000001100000,
31'b0000000000001000000001010000100,
31'b0001000000100000010001000000000,
31'b0000000000000000100000101000000,
31'b0001000010000000000000001100000,
31'b0000000000000000000001010000100,
31'b1000000010000000110000000000100,
31'b0000000000001000100000101000000,
31'b0101000111000000000000000000000,
31'b1000010000000000100100001000000,
31'b0001001000000000000000000000110,
31'b1000100000000000001100000000100,
31'b1000000000000010001000010010000,
31'b1000000000000000001000010010000,
31'b0010100000000001000000001000100,
31'b1100100000000000000000101000000,
31'b0100000000000000010010000000010,
31'b0110000100000000000000000101000,
31'b0100001100000000000000100000000,
31'b0100010000000000010000001001000,
31'b0100000100000000101000000010000,
31'b0010000000000000001000000000110,
31'b1100000000000000010000000010001,
31'b0010010010000001000000000001000,
31'b1010010000000000000000000010001,
31'b0010000000001000000000001001000,
31'b0011000001000000000000001010000,
31'b0010000001000000000011000000001,
31'b0010000000000010000000001001000,
31'b0010000000000000000000001001000,
31'b0010010000000000000010000000010,
31'b0010000000000100000000001001000,
31'b1100000100000001000000000000001,
31'b0010000100000000000000100000101,
31'b0100001100100000000000100000000,
31'b0000000100000001000001000001000,
31'b0010110010000000000000000000100,
31'b0010000000010000000000001001000,
31'b1100000000000000100010100000000,
31'b0010000000010100000000001001000,
31'b0101001000000000000000000000000,
31'b0101001000000010000000000000000,
31'b0101001000000100000000000000000,
31'b0110000000011000001000000000000,
31'b0101001000001000000000000000000,
31'b0110000000010100001000000000000,
31'b0110000000010010001000000000000,
31'b0110000000010000001000000000000,
31'b0101001000010000000000000000000,
31'b0110000000001100001000000000000,
31'b0000000000000000010010000000100,
31'b0110000000001000001000000000000,
31'b0110000000000110001000000000000,
31'b0110000000000100001000000000000,
31'b0110000000000010001000000000000,
31'b0110000000000000001000000000000,
31'b0101001000100000000000000000000,
31'b0000010000000000011000000000000,
31'b0101001000100100000000000000000,
31'b0011000000000000000000000000101,
31'b0110010000000000000010000000100,
31'b0001000000010000000010010000000,
31'b1000100010000000100000100000000,
31'b0110000000110000001000000000000,
31'b0101001000110000000000000000000,
31'b0001000000001000000010010000000,
31'b0100010000000000000000010000001,
31'b0110000000101000001000000000000,
31'b0001000000000010000010010000000,
31'b0001000000000000000010010000000,
31'b0110000000100010001000000000000,
31'b0110000000100000001000000000000,
31'b0101001001000000000000000000000,
31'b0101001001000010000000000000000,
31'b0100000010010000000000100000000,
31'b0100001000001000000000000011000,
31'b1001000100000000000000010100000,
31'b1001001000000000000010001000000,
31'b0100001000000010000000000011000,
31'b0100001000000000000000000011000,
31'b0100000010000100000000100000000,
31'b0101000000001000100000000100000,
31'b0100000010000000000000100000000,
31'b0100000010000010000000100000000,
31'b0101000000000010100000000100000,
31'b0101000000000000100000000100000,
31'b0100000010001000000000100000000,
31'b0000000000000001000110000000000,
31'b0101001001100000000000000000000,
31'b0001000100000000100000001000000,
31'b0100001000000001000100010000000,
31'b1010100000000000101000000000000,
31'b0010010010000000010000100000000,
31'b0001000100001000100000001000000,
31'b0000000010000000000100000001010,
31'b0100001000100000000000000011000,
31'b1101000000000000000000011000000,
31'b0001000100010000100000001000000,
31'b0100000010100000000000100000000,
31'b0100000010100010000000100000000,
31'b1001101000000000100000000000000,
31'b0001000001000000000010010000000,
31'b0100000010101000000000100000000,
31'b0100000000000000000001010000010,
31'b0000100000000000010000000000010,
31'b0100000000000000001000000110000,
31'b0100000001010000000000100000000,
31'b0100000001010010000000100000000,
31'b0110000000000000100000000001000,
31'b0110000000000010100000000001000,
31'b1010000000010000010100000000000,
31'b1010000000000000100001000000001,
31'b0100000001000100000000100000000,
31'b0100000001000110000000100000000,
31'b0100000001000000000000100000000,
31'b0100000001000010000000100000000,
31'b1010000000000100010100000000000,
31'b1010000100000000000000010001000,
31'b1010000000000000010100000000000,
31'b1000000000000000000010101000000,
31'b1100010000000000000100000000000,
31'b0001000000000000000100000010010,
31'b1100010000000100000100000000000,
31'b0011000010000000000000000000101,
31'b1100010000001000000100000000000,
31'b0001000010010000000010010000000,
31'b1000100000000000100000100000000,
31'b1001000000000000000110000000001,
31'b1100010000010000000100000000000,
31'b0001000010001000000010010000000,
31'b0100000001100000000000100000000,
31'b0100010100000000001001000000000,
31'b0001001000000001000001000010000,
31'b0001000010000000000010010000000,
31'b1010000000100000010100000000000,
31'b1011100000000000000000000010000,
31'b0100000000010100000000100000000,
31'b0100000001000000001000000110000,
31'b0100000000010000000000100000000,
31'b0100000000010010000000100000000,
31'b0110000001000000100000000001000,
31'b1000000100000000000001001000100,
31'b0100000000011000000000100000000,
31'b0100001010000000000000000011000,
31'b0100000000000100000000100000000,
31'b0100000000000110000000100000000,
31'b0100000000000000000000100000000,
31'b0100000000000010000000100000000,
31'b0100000000001100000000100000000,
31'b0101000010000000100000000100000,
31'b0100000000001000000000100000000,
31'b0100000000001010000000100000000,
31'b1100010001000000000100000000000,
31'b0001000110000000100000001000000,
31'b0100000000110000000000100000000,
31'b0100000000110010000000100000000,
31'b0010010000000000010000100000000,
31'b0000010000000000000110001000000,
31'b0000000000000000000100000001010,
31'b0000001000000000000010110000000,
31'b1010100000000000000000000001000,
31'b1100000000000000000001000100100,
31'b0100000000100000000000100000000,
31'b0100000000100010000000100000000,
31'b1100000000000000110000000000010,
31'b0001010000000000110000000010000,
31'b0100000000101000000000100000000,
31'b0100000010000000000001010000010,
31'b0101001100000000000000000000000,
31'b0101001100000010000000000000000,
31'b0101001100000100000000000000000,
31'b1000010000100000100000000000001,
31'b1110000000000000000101000000000,
31'b0010000010000000011001000000000,
31'b1010000000000000101000010000000,
31'b0010000000000000000100000001001,
31'b0001100001000000000010000000000,
31'b1001001000000000100000010000000,
31'b0100100000000000000001000000010,
31'b0110000100001000001000000000000,
31'b0001100001001000000010000000000,
31'b1101100000000000000000001000000,
31'b0110000100000010001000000000000,
31'b0110000100000000001000000000000,
31'b0101001100100000000000000000000,
31'b0001000001000000100000001000000,
31'b1000010000000010100000000000001,
31'b1000010000000000100000000000001,
31'b1101000000000000100010000000000,
31'b0001000100010000000010010000000,
31'b1000000000000001000100000100000,
31'b1000010000001000100000000000001,
31'b0010100000000001000000000100010,
31'b0001000100001000000010010000000,
31'b1000010000000000010101000000000,
31'b1000010000010000100000000000001,
31'b0001001000000000000000001100000,
31'b0001000100000000000010010000000,
31'b1000001000000000110000000000100,
31'b0110000100100000001000000000000,
31'b0000000000000000010001100000000,
31'b0001000000100000100000001000000,
31'b0001000010000000000000000000110,
31'b1000000010000000100000110000000,
31'b1001000000000000000000010100000,
31'b1001000000000010000000010100000,
31'b1001000000000100000000010100000,
31'b0100110000010000000000000000001,
31'b0001100000000000000010000000000,
31'b0001100000000010000010000000000,
31'b0100000110000000000000100000000,
31'b0100110000001000000000000000001,
31'b0001100000001000000010000000000,
31'b0101000100000000100000000100000,
31'b0100110000000010000000000000001,
31'b0100110000000000000000000000001,
31'b0001000000000010100000001000000,
31'b0001000000000000100000001000000,
31'b1000000000001000100001000000010,
31'b1000000000000000010000000100100,
31'b1001000000100000000000010100000,
31'b0001000000001000100000001000000,
31'b1000000000000000100001000000010,
31'b1000000000001000010000000100100,
31'b0010000000000000000000101010000,
31'b0001000000010000100000001000000,
31'b0110100000000000001000010000000,
31'b1000001000000001100100000000000,
31'b0010111000000000000000000000100,
31'b0001000101000000000010010000000,
31'b1000011000000000000000000100001,
31'b1000010000000001000001000000100,
31'b0100000000000000000011000000100,
31'b0100000100000000001000000110000,
31'b0001000001000000000000000000110,
31'b1000000001000000100000110000000,
31'b0110000100000000100000000001000,
31'b0010000000000000011001000000000,
31'b0001011000000001000000000100000,
31'b0010000010000000000100000001001,
31'b0100000101000100000000100000000,
31'b1010000000001000000000010001000,
31'b0100000101000000000000100000000,
31'b0100010000100000001001000000000,
31'b1010000000000010000000010001000,
31'b1010000000000000000000010001000,
31'b1010000100000000010100000000000,
31'b1010000000000100000000010001000,
31'b1100010100000000000100000000000,
31'b0001000100000000000100000010010,
31'b0011001000000000000000001010000,
31'b1100000000000000000010100100000,
31'b0000100000000101000000000010010,
31'b0000000001000000010000010000010,
31'b0000100000000001000000000010010,
31'b0100100000010000000000110000000,
31'b1010000000000001000100000010000,
31'b0000010000000000100100010000000,
31'b0100010000000010001001000000000,
31'b0100010000000000001001000000000,
31'b0000000000000010001000001010000,
31'b0000000000000000001000001010000,
31'b0100100000000010000000110000000,
31'b0100100000000000000000110000000,
31'b0001000000000100000000000000110,
31'b1000000000001000000001001000100,
31'b0001000000000000000000000000110,
31'b1000000000000000100000110000000,
31'b1001000010000000000000010100000,
31'b1000000000000000000001001000100,
31'b0001000000001000000000000000110,
31'b1000000000001000100000110000000,
31'b0100000100000100000000100000000,
31'b0100010000000000000110000100000,
31'b0100000100000000000000100000000,
31'b0100000100000010000000100000000,
31'b0100000100001100000000100000000,
31'b1010000001000000000000010001000,
31'b0100000100001000000000100000000,
31'b0100110010000000000000000000001,
31'b0001000010000010100000001000000,
31'b0001000010000000100000001000000,
31'b0001000000100000000000000000110,
31'b1000000010000000010000000100100,
31'b0000000000000100000000101100000,
31'b0000000000000000010000010000010,
31'b0000000000000000000000101100000,
31'b0000000000000100010000010000010,
31'b1100000000000000001010000010000,
31'b0001010000000000001010000000010,
31'b0100000100100000000000100000000,
31'b0100010001000000001001000000000,
31'b0100000000000100001000000000011,
31'b0000000001000000001000001010000,
31'b0100000000000000001000000000011,
31'b0100100001000000000000110000000,
31'b0101010000000000000000000000000,
31'b1000000000000000000000000010010,
31'b0101010000000100000000000000000,
31'b0000000000001000000010000000001,
31'b0101010000001000000000000000000,
31'b0000000000000100000010000000001,
31'b0000000000000010000010000000001,
31'b0000000000000000000010000000001,
31'b0101010000010000000000000000000,
31'b0010000000000000000000010000100,
31'b0101010000010100000000000000000,
31'b0010000000000100000000010000100,
31'b0101010000011000000000000000000,
31'b0010000000001000000000010000100,
31'b0011000000100000010000000000000,
31'b0000000000010000000010000000001,
31'b0101010000100000000000000000000,
31'b0000001000000000011000000000000,
31'b0101010000100100000000000000000,
31'b0000001000000100011000000000000,
31'b0110001000000000000010000000100,
31'b0000001000001000011000000000000,
31'b0011000000010000010000000000000,
31'b0000000000100000000010000000001,
31'b0101010000110000000000000000000,
31'b0010000000100000000000010000100,
31'b0100001000000000000000010000001,
31'b0101000000000000001010000000100,
31'b0011000000000100010000000000000,
31'b0011000000000110010000000000000,
31'b0011000000000000010000000000000,
31'b0011000000000010010000000000000,
31'b0101010001000000000000000000000,
31'b0000000000000000000001001001000,
31'b1100000000000000000000001000001,
31'b0000000001001000000010000000001,
31'b1001000000000100000000000001010,
31'b0000000001000100000010000000001,
31'b1001000000000000000000000001010,
31'b0000000001000000000010000000001,
31'b0101010001010000000000000000000,
31'b0010000001000000000000010000100,
31'b1100000000010000000000001000001,
31'b0010000100001001000000000001000,
31'b0010100100100000000000000000100,
31'b0010000100000101000000000001000,
31'b1001000000010000000000000001010,
31'b0010000100000001000000000001000,
31'b0101010001100000000000000000000,
31'b0000001001000000011000000000000,
31'b1100000000100000000000001000001,
31'b0000101000000000000000001100001,
31'b0010100100010000000000000000100,
31'b0000001010000000000110001000000,
31'b1001000000100000000000000001010,
31'b0000000010000000010000000101000,
31'b0010100100001000000000000000100,
31'b0010000000000000010000000011000,
31'b1101000000000000000100100000000,
31'b0011000000000001000100000000100,
31'b0010100100000000000000000000100,
31'b0100100000000000100000000010010,
31'b1000000100000000000000000100001,
31'b1001000010000001000010000000000,
31'b0101010010000000000000000000000,
31'b0000100000000000000100000100000,
31'b0101010010000100000000000000000,
31'b0000100000000100000100000100000,
31'b0101010010001000000000000000000,
31'b0000100000001000000100000100000,
31'b0001000100000001000000000100000,
31'b0000000010000000000010000000001,
31'b0101010010010000000000000000000,
31'b0010000010000000000000010000100,
31'b0101000000100001000000001000000,
31'b1010000000001000000000000100010,
31'b1000001000000000000000100001010,
31'b1000000000000000000110010000000,
31'b1010000000000010000000000100010,
31'b1010000000000000000000000100010,
31'b1100001000000000000100000000000,
31'b0000100000100000000100000100000,
31'b1100001000000100000100000000000,
31'b0000100001000000001011000000000,
31'b1100001000001000000100000000000,
31'b0000100000101000000100000100000,
31'b0011000010010000010000000000000,
31'b0000000010100000000010000000001,
31'b1100001000010000000100000000000,
31'b0010000010100000000000010000100,
31'b0101000000000001000000001000000,
31'b0101000000000011000000001000000,
31'b0011000010000100010000000000000,
31'b1100000000000001000001000000010,
31'b0011000010000000010000000000000,
31'b1010000000100000000000000100010,
31'b0101010011000000000000000000000,
31'b0000100001000000000100000100000,
31'b1100000010000000000000001000001,
31'b0000100001000100000100000100000,
31'b0010001000100000010000100000000,
31'b0000101000000000010001000000001,
31'b1010000000000001010000000000001,
31'b0000000011000000000010000000001,
31'b0100000000000000000100011000000,
31'b0110010000000000000000000101000,
31'b0100011000000000000000100000000,
31'b0100011000000010000000100000000,
31'b0000101000000000100100000000000,
31'b1001000000000000101000000000010,
31'b0100100000000000000000001010100,
31'b1010000001000000000000000100010,
31'b1100001001000000000100000000000,
31'b0000100001100000000100000100000,
31'b0010000100001000000010000000010,
31'b0000100000000000001011000000000,
31'b0010001000000000010000100000000,
31'b0000001000000000000110001000000,
31'b0010000100000000000010000000010,
31'b0000000000000000010000000101000,
31'b1100010000000001000000000000001,
31'b0010010000000000000000100000101,
31'b0101000001000001000000001000000,
31'b0001000000000000011000100000000,
31'b0010100110000000000000000000100,
31'b1100000000000000100100000100000,
31'b1001000000000011000010000000000,
31'b1001000000000001000010000000000,
31'b0101010100000000000000000000000,
31'b0000000000000001100000100000000,
31'b0101010100000100000000000000000,
31'b0000000100001000000010000000001,
31'b0101010100001000000000000000000,
31'b0000000100000100000010000000001,
31'b0001000010000001000000000100000,
31'b0000000100000000000010000000001,
31'b0011000000000001000000000010000,
31'b0010000100000000000000010000100,
31'b0011000000000101000000000010000,
31'b0010000100000100000000010000100,
31'b0011000000001001000000000010000,
31'b0010000100001000000000010000100,
31'b1000000010000000010010000001000,
31'b0010000001000001000000000001000,
31'b0101010100100000000000000000000,
31'b0000001100000000011000000000000,
31'b1000001000000010100000000000001,
31'b1000001000000000100000000000001,
31'b0111000010000000000001000000000,
31'b1000000000000101010000000000010,
31'b1000000001010000000000000100001,
31'b1000000000000001010000000000010,
31'b0011000000100001000000000010000,
31'b0010100000000001010100000000000,
31'b1000001000000000010101000000000,
31'b1000010000000000000001000100010,
31'b0010100001000000000000000000100,
31'b0100100010000000000100001000000,
31'b1000000001000000000000000100001,
31'b1000000001000010000000000100001,
31'b0101010101000000000000000000000,
31'b0000000100000000000001001001000,
31'b1100000100000000000000001000001,
31'b0010000000011001000000000001000,
31'b0010100000110000000000000000100,
31'b0010000000010101000000000001000,
31'b1001000100000000000000000001010,
31'b0010000000010001000000000001000,
31'b0011000001000001000000000010000,
31'b0010000101000000000000010000100,
31'b1000000000101000000000000100001,
31'b0010000000001001000000000001000,
31'b0010100000100000000000000000100,
31'b0010000000000101000000000001000,
31'b1000000000100000000000000100001,
31'b0010000000000001000000000001000,
31'b1010000010000000000000000010001,
31'b0101000000000000001001100000000,
31'b1000000000000000000100000000110,
31'b1000001001000000100000000000001,
31'b0010100000010000000000000000100,
31'b0101110000000000000000010000000,
31'b1000000000010000000000000100001,
31'b1000000001000001010000000000010,
31'b0010100000001000000000000000100,
31'b0100100000000000011010000000000,
31'b1000000000001000000000000100001,
31'b1000010000000001100100000000000,
31'b0010100000000000000000000000100,
31'b0100000000000000000001000101000,
31'b1000000000000000000000000100001,
31'b1000000000000010000000000100001,
31'b0101010110000000000000000000000,
31'b0000100100000000000100000100000,
31'b0001000000001001000000000100000,
31'b0001010000000000100100000000001,
31'b0100000000000000100110000000000,
31'b0101100000000000000000100000001,
31'b0001000000000001000000000100000,
31'b0001000000000011000000000100000,
31'b0011000010000001000000000010000,
31'b0010001000000001001000000100000,
31'b0001010000000000010001000000000,
31'b0100001000100000001001000000000,
31'b1000001000000000000100001100000,
31'b1000010000000000010000001000010,
31'b1000000000000000010010000001000,
31'b1010000100000000000000000100010,
31'b1100001100000000000100000000000,
31'b0000100100100000000100000100000,
31'b0011010000000000000000001010000,
31'b1110000000000000000000001000010,
31'b0111000000000000000001000000000,
31'b0111000000000010000001000000000,
31'b0010000001000000000010000000010,
31'b1011000000000000000000000001001,
31'b1000100001000000000110000000000,
31'b0000100000000000001000100000100,
31'b0101000100000001000000001000000,
31'b0100001000000000001001000000000,
31'b0111000000010000000001000000000,
31'b0100100000000000000100001000000,
31'b1000000011000000000000000100001,
31'b0100100000000100000100001000000,
31'b1010000000100000000000000010001,
31'b1000000000000000100100001000000,
31'b0010001000000001000000100010000,
31'b1100001000000000000000000010100,
31'b0010000000000001101000000000000,
31'b1000010000000000001000010010000,
31'b0010000000100000000010000000010,
31'b0010000010010001000000000001000,
31'b1000100000100000000110000000000,
31'b1001000000000000010010000010000,
31'b0100011100000000000000100000000,
31'b0100000000000000010000001001000,
31'b0010100010100000000000000000100,
31'b0010010000000000001000000000110,
31'b1000000010100000000000000100001,
31'b0010000010000001000000000001000,
31'b1010000000000000000000000010001,
31'b1010000000000010000000000010001,
31'b0010000000001000000010000000010,
31'b0110000000000000000001000011000,
31'b0000000000000000000100010100000,
31'b0010010000000000000000001001000,
31'b0010000000000000000010000000010,
31'b0010000000000010000010000000010,
31'b1000100000000000000110000000000,
31'b1001000000000000100000100000001,
31'b1000100000000100000110000000000,
31'b0100001001000000001001000000000,
31'b0010100010000000000000000000100,
31'b0100100001000000000100001000000,
31'b1000000010000000000000000100001,
31'b1001000100000001000010000000000,
31'b0101011000000000000000000000000,
31'b0000000000100000011000000000000,
31'b0101011000000100000000000000000,
31'b0000001000001000000010000000001,
31'b0110000000100000000010000000100,
31'b0000001000000100000010000000001,
31'b0001000000000000001000010000100,
31'b0000001000000000000010000000001,
31'b0101011000010000000000000000000,
31'b0010001000000000000000010000100,
31'b0100000000100000000000010000001,
31'b0110010000001000001000000000000,
31'b1000000010000000000000100001010,
31'b0110010000000100001000000000000,
31'b0110010000000010001000000000000,
31'b0110010000000000001000000000000,
31'b0000000000000010011000000000000,
31'b0000000000000000011000000000000,
31'b0100000000010000000000010000001,
31'b0000000000000100011000000000000,
31'b0110000000000000000010000000100,
31'b0000000000001000011000000000000,
31'b0110000000000100000010000000100,
31'b0000001000100000000010000000001,
31'b0100000000000100000000010000001,
31'b0000000000010000011000000000000,
31'b0100000000000000000000010000001,
31'b0100000000000010000000010000001,
31'b0110000000010000000010000000100,
31'b0001010000000000000010010000000,
31'b0100000000001000000000010000001,
31'b0110010000100000001000000000000,
31'b0101011001000000000000000000000,
31'b0000001000000000000001001001000,
31'b1100001000000000000000001000001,
31'b0000100000100000000000001100001,
31'b0010000010100000010000100000000,
31'b0000100010000000010001000000001,
31'b1001001000000000000000000001010,
31'b0000100000000000001100000001000,
31'b0101000000000001000100000000001,
31'b1010000000000000001000000001010,
31'b0100010010000000000000100000000,
31'b0100100100001000000000000000001,
31'b0000100010000000100100000000000,
31'b0101010000000000100000000100000,
31'b0100100100000010000000000000001,
31'b0100100100000000000000000000001,
31'b0100000000000001000000101000000,
31'b0000000001000000011000000000000,
31'b0100000001010000000000010000001,
31'b0000100000000000000000001100001,
31'b0010000010000000010000100000000,
31'b0000000010000000000110001000000,
31'b0011000000000000000001000000110,
31'b0000100000100000001100000001000,
31'b0100000001000100000000010000001,
31'b0000000001010000011000000000000,
31'b0100000001000000000000010000001,
31'b0100100000000000001000100000010,
31'b0010101100000000000000000000100,
31'b0001010001000000000010010000000,
31'b1001000000000000000001010010000,
31'b1000000100000001000001000000100,
31'b1100000000100000000100000000000,
31'b0000101000000000000100000100000,
31'b1100000000100100000100000000000,
31'b0000101000000100000100000100000,
31'b1100000000101000000100000000000,
31'b0000101000001000000100000100000,
31'b0001001100000001000000000100000,
31'b0000001010000000000010000000001,
31'b1100000000110000000100000000000,
31'b0010001010000000000000010000100,
31'b0100010001000000000000100000000,
31'b0100010001000010000000100000000,
31'b1000000000000000000000100001010,
31'b1000001000000000000110010000000,
31'b1010010000000000010100000000000,
31'b1010001000000000000000000100010,
31'b1100000000000000000100000000000,
31'b0000000010000000011000000000000,
31'b1100000000000100000100000000000,
31'b0000000010000100011000000000000,
31'b1100000000001000000100000000000,
31'b0000000010001000011000000000000,
31'b1100000000001100000100000000000,
31'b0000001010100000000010000000001,
31'b1100000000010000000100000000000,
31'b0000000100000000100100010000000,
31'b0000000000000000110000000001000,
31'b0100000100000000001001000000000,
31'b1100000000011000000100000000000,
31'b0001010010000000000010010000000,
31'b0110100000000000000000000000010,
31'b0110100000000010000000000000010,
31'b1100000001100000000100000000000,
31'b0000101001000000000100000100000,
31'b1010000000000000100000000000010,
31'b1100000100000000000000000010100,
31'b0010000000100000010000100000000,
31'b0000100000000000010001000000001,
31'b1100100000000000010000000001000,
31'b0000100010000000001100000001000,
31'b0100010000000100000000100000000,
31'b0100010000000110000000100000000,
31'b0100010000000000000000100000000,
31'b0100010000000010000000100000000,
31'b0000100000000000100100000000000,
31'b0001000000000000000010100000001,
31'b0100010000001000000000100000000,
31'b0100100110000000000000000000001,
31'b1100000001000000000100000000000,
31'b0000000011000000011000000000000,
31'b1100000001000100000100000000000,
31'b0000101000000000001011000000000,
31'b0010000000000000010000100000000,
31'b0000000000000000000110001000000,
31'b0010000000000100010000100000000,
31'b0000001000000000010000000101000,
31'b1100000001010000000100000000000,
31'b0001000100000000001010000000010,
31'b0100010000100000000000100000000,
31'b0100010000100010000000100000000,
31'b0010000000010000010000100000000,
31'b0001000000000000110000000010000,
31'b0110100001000000000000000000010,
31'b1001001000000001000010000000000,
31'b0101011100000000000000000000000,
31'b0000001000000001100000100000000,
31'b1010000000000000000100001010000,
31'b1000000000100000100000000000001,
31'b0000100001000000011000010000000,
31'b0000000000000101001000000010000,
31'b0000000000000011001000000010000,
31'b0000000000000001001000000010000,
31'b0011001000000001000000000010000,
31'b0010001100000000000000010000100,
31'b1000100000000000000010001000001,
31'b1001100000000000000001000010000,
31'b0000100000000000000000001010010,
31'b0100100001000100000000000000001,
31'b0100100001000010000000000000001,
31'b0100100001000000000000000000001,
31'b0100000000000000100001000001000,
31'b0000000100000000011000000000000,
31'b1000000000000010100000000000001,
31'b1000000000000000100000000000001,
31'b0110000100000000000010000000100,
31'b0000000100001000011000000000000,
31'b1000010000000001000100000100000,
31'b1000000000001000100000000000001,
31'b1000000010000000001000000001001,
31'b0000000100010000011000000000000,
31'b1000000000000000010101000000000,
31'b1000000000010000100000000000001,
31'b0011000000000000000010100000010,
31'b0001010100000000000010010000000,
31'b1000001001000000000000000100001,
31'b1000000001000001000001000000100,
31'b0001000000000001001000000001000,
31'b0001010000100000100000001000000,
31'b0010000010000001000000100010000,
31'b1100000010000000000000000010100,
31'b0000100000000000011000010000000,
31'b0100100000010100000000000000001,
31'b0100100000010010000000000000001,
31'b0100100000010000000000000000001,
31'b0001110000000000000010000000000,
31'b0100100000001100000000000000001,
31'b0100100000001010000000000000001,
31'b0100100000001000000000000000001,
31'b0000000000000001000000100100000,
31'b0100100000000100000000000000001,
31'b0100100000000010000000000000001,
31'b0100100000000000000000000000001,
31'b0100000100000001000000101000000,
31'b0001010000000000100000001000000,
31'b1000001000000000000100000000110,
31'b1000000001000000100000000000001,
31'b0010101000010000000000000000100,
31'b0001010000001000100000001000000,
31'b1000010000000000100001000000010,
31'b1000000001001000100000000000001,
31'b0010101000001000000000000000100,
31'b0001010000010000100000001000000,
31'b1000001000001000000000000100001,
31'b1000000001010000100000000000001,
31'b0010101000000000000000000000100,
31'b1010000000000000000000100001001,
31'b1000001000000000000000000100001,
31'b1000000000000001000001000000100,
31'b1100000100100000000100000000000,
31'b0010100000000000010000110000000,
31'b0010100000000000000000001100010,
31'b1100000001000000000000000010100,
31'b1101000000000000000000000001100,
31'b0011000000000001000000100001000,
31'b0001001000000001000000000100000,
31'b0001000000000000000001000000101,
31'b1000000000100000001000000001001,
31'b0010000000000001001000000100000,
31'b0100010101000000000000100000000,
31'b0100000000100000001001000000000,
31'b1000000000000000000100001100000,
31'b1010010000000000000000010001000,
31'b1000001000000000010010000001000,
31'b0100100011000000000000000000001,
31'b1100000100000000000100000000000,
31'b0000000110000000011000000000000,
31'b1100000100000100000100000000000,
31'b1000000010000000100000000000001,
31'b1100000100001000000100000000000,
31'b0000010001000000010000010000010,
31'b0011100000000000000000100000100,
31'b1101100000000001000000000000000,
31'b1000000000000000001000000001001,
31'b0000000000000000100100010000000,
31'b0100000000000010001001000000000,
31'b0100000000000000001001000000000,
31'b1000000000100000000100001100000,
31'b0000010000000000001000001010000,
31'b0110100100000000000000000000010,
31'b0100000000001000001001000000000,
31'b0010000000000101000000100010000,
31'b1100000000000100000000000010100,
31'b0010000000000001000000100010000,
31'b1100000000000000000000000010100,
31'b0010001000000001101000000000000,
31'b1100100000000000000100010000000,
31'b0010001000100000000010000000010,
31'b1100000000001000000000000010100,
31'b0100010100000100000000100000000,
31'b0100000000000000000110000100000,
31'b0100010100000000000000100000000,
31'b0001000000000001100000000000000,
31'b0000100100000000100100000000000,
31'b0100100010000100000000000000001,
31'b0100100010000010000000000000001,
31'b0100100010000000000000000000001,
31'b1100000101000000000100000000000,
31'b0001010010000000100000001000000,
31'b0010001000001000000010000000010,
31'b1100000000100000000000000010100,
31'b0010000100000000010000100000000,
31'b0000010000000000010000010000010,
31'b0010001000000000000010000000010,
31'b0010001000000010000010000000010,
31'b1000101000000000000110000000000,
31'b0001000000000000001010000000010,
31'b0100010100100000000000100000000,
31'b0100000001000000001001000000000,
31'b0010101010000000000000000000100,
31'b0001000100000000110000000010000,
31'b1000001010000000000000000100001,
31'b1001000000000000001000000010001,
31'b0101100000000000000000000000000,
31'b0101100000000010000000000000000,
31'b0101100000000100000000000000000,
31'b0101100000000110000000000000000,
31'b0101100000001000000000000000000,
31'b0101100000001010000000000000000,
31'b0101100000001100000000000000000,
31'b0100000100000001000100000000000,
31'b0101100000010000000000000000000,
31'b0110000000000000000101001000000,
31'b0101100000010100000000000000000,
31'b1000010000000000000000010100001,
31'b1100000000000001001001000000000,
31'b0010010000000100000100000010000,
31'b1010000000100000001000000100000,
31'b0010010000000000000100000010000,
31'b1000000010000000001000000010000,
31'b1001001000000000000000000100000,
31'b1011000000000000000000100001000,
31'b1001001000000100000000000100000,
31'b1001000001010000100000000000000,
31'b1010000001000000000000100010000,
31'b1010000000010000001000000100000,
31'b0100100000000000010000010000100,
31'b1001000001001000100000000000000,
31'b1001001000010000000000000100000,
31'b1010000000001000001000000100000,
31'b1000000000000000100000000011000,
31'b1001000001000000100000000000000,
31'b1001000001000010100000000000000,
31'b1010000000000000001000000100000,
31'b1010000000000010001000000100000,
31'b0101100001000000000000000000000,
31'b0101100001000010000000000000000,
31'b0100000100000000010000000000100,
31'b0100100000001000000000000011000,
31'b1001000000110000100000000000000,
31'b1010000000100000000000100010000,
31'b0100100000000010000000000011000,
31'b0100100000000000000000000011000,
31'b0000000010000000000001000000100,
31'b0001000000000000000000011100000,
31'b0001000000000000010000100000010,
31'b1000000010100000000000100100000,
31'b1001000000100000100000000000000,
31'b1001000000100010100000000000000,
31'b1001000000100100100000000000000,
31'b0100100000010000000000000011000,
31'b1001000000011000100000000000000,
31'b1010000000001000000000100010000,
31'b0100100000000001000100010000000,
31'b1010001000000000101000000000000,
31'b1001000000010000100000000000000,
31'b1010000000000000000000100010000,
31'b1001000000010100100000000000000,
31'b1010000000000100000000100010000,
31'b1001000000001000100000000000000,
31'b1001000000001010100000000000000,
31'b1001000000001100100000000000000,
31'b1000000010000000000000100100000,
31'b1001000000000000100000000000000,
31'b1001000000000010100000000000000,
31'b1001000000000100100000000000000,
31'b1001000000000110100000000000000,
31'b0000001000000000010000000000010,
31'b0000010000000000000100000100000,
31'b0000000100000000000010100000000,
31'b0000010000000100000100000100000,
31'b0000000000000001100000000000001,
31'b0000010000001000000100000100000,
31'b0000000100001000000010100000000,
31'b0100100000000000100000100100000,
31'b0000000001000000000001000000100,
31'b0000010000010000000100000100000,
31'b0000000100010000000010100000000,
31'b1000010000000000000010000010100,
31'b0000000001001000000001000000100,
31'b0000010000000000000000000000111,
31'b0000000100011000000010100000000,
31'b0011000000000000011000000000010,
31'b1000000000000000001000000010000,
31'b1000000000000010001000000010000,
31'b1000000000000100001000000010000,
31'b1000000001010000000000100100000,
31'b1000000000001000001000000010000,
31'b1010000000000000100000000101000,
31'b1000001000000000100000100000000,
31'b1001000001000000001000000001000,
31'b1000000000010000001000000010000,
31'b1000000001000100000000100100000,
31'b1000000001000010000000100100000,
31'b1000000001000000000000100100000,
31'b1001000011000000100000000000000,
31'b0100010100000000000100001000000,
31'b1010000010000000001000000100000,
31'b1011001000000000000000000010000,
31'b0000000000010000000001000000100,
31'b0000010001000000000100000100000,
31'b0000000101000000000010100000000,
31'b1000000100000000001100000000100,
31'b0000000001000001100000000000001,
31'b0000011000000000010001000000001,
31'b0010000100000001000000001000100,
31'b1100000100000000000000101000000,
31'b0000000000000000000001000000100,
31'b0000000000000010000001000000100,
31'b0000000000000100000001000000100,
31'b1000000000100000000000100100000,
31'b0000000000001000000001000000100,
31'b0000000000001010000001000000100,
31'b0000000000001100000001000000100,
31'b1001000000000000000000001000110,
31'b1000000001000000001000000010000,
31'b1000000001000010001000000010000,
31'b1000000001000100001000000010000,
31'b1000000000010000000000100100000,
31'b1001000010010000100000000000000,
31'b1010000010000000000000100010000,
31'b1001000000000010001000000001000,
31'b1001000000000000001000000001000,
31'b0000000000100000000001000000100,
31'b1000000000000100000000100100000,
31'b1000000000000010000000100100000,
31'b1000000000000000000000100100000,
31'b1001000010000000100000000000000,
31'b1001000010000010100000000000000,
31'b1001000010000100100000000000000,
31'b1000000000001000000000100100000,
31'b0101100100000000000000000000000,
31'b0101100100000010000000000000000,
31'b0000000010000000000010100000000,
31'b0100000000001001000100000000000,
31'b0101100100001000000000000000000,
31'b0100000000000101000100000000000,
31'b0100000000000011000100000000000,
31'b0100000000000001000100000000000,
31'b0001001001000000000010000000000,
31'b1001100000000000100000010000000,
31'b0100001000000000000001000000010,
31'b0100001000000010000001000000010,
31'b0010010001100000000000000000100,
31'b1101001000000000000000001000000,
31'b0100001000001000000001000000010,
31'b0100000000010001000100000000000,
31'b1001000000000000000010011000000,
31'b1001001100000000000000000100000,
31'b0100000000000000000000010011000,
31'b0100000000101001000100000000000,
31'b0101000001000010000000010000000,
31'b0101000001000000000000010000000,
31'b0100000000100011000100000000000,
31'b0100000000100001000100000000000,
31'b0010010001001000000000000000100,
31'b0010010000000001010100000000000,
31'b0100001000100000000001000000010,
31'b0000000010000000000101000010000,
31'b0010010001000000000000000000100,
31'b0101000001010000000000010000000,
31'b1010000100000000001000000100000,
31'b0100001010000000000000110000000,
31'b0100000000000100010000000000100,
31'b0101000000101000000000010000000,
31'b0100000000000000010000000000100,
31'b0100000000000010010000000000100,
31'b0101000000100010000000010000000,
31'b0101000000100000000000010000000,
31'b0100000000001000010000000000100,
31'b0010000000000000001010000000000,
31'b0001001000000000000010000000000,
31'b0001001000000010000010000000000,
31'b0100000000010000010000000000100,
31'b0100011000001000000000000000001,
31'b0010010000100000000000000000100,
31'b0101000000110000000000010000000,
31'b0100011000000010000000000000001,
31'b0100011000000000000000000000001,
31'b0101000000001010000000010000000,
31'b0101000000001000000000010000000,
31'b0100000000100000010000000000100,
31'b0101000000001100000000010000000,
31'b0101000000000010000000010000000,
31'b0101000000000000000000010000000,
31'b0101000000000110000000010000000,
31'b0101000000000100000000010000000,
31'b0010010000001000000000000000100,
31'b0101000000011000000000010000000,
31'b0110001000000000001000010000000,
31'b1000100000000001100100000000000,
31'b0010010000000000000000000000100,
31'b0101000000010000000000010000000,
31'b0010010000000100000000000000100,
31'b0101000000010100000000010000000,
31'b0000000000000100000010100000000,
31'b0000010100000000000100000100000,
31'b0000000000000000000010100000000,
31'b0000000000000010000010100000000,
31'b0000000100000001100000000000001,
31'b0101010000000000000000100000001,
31'b0000000000001000000010100000000,
31'b0100000010000001000100000000000,
31'b0000000101000000000001000000100,
31'b0000010100010000000100000100000,
31'b0000000000010000000010100000000,
31'b0000000000100000000101000010000,
31'b0010000001000000100010000001000,
31'b1100000000000001000000010000001,
31'b0000000000011000000010100000000,
31'b0100001000100000000000110000000,
31'b1000000100000000001000000010000,
31'b1000000100000010001000000010000,
31'b0000000000100000000010100000000,
31'b0000000000100010000010100000000,
31'b1000000100001000001000000010000,
31'b0101000011000000000000010000000,
31'b0000001000000001000000000010010,
31'b0100001000010000000000110000000,
31'b1000010001000000000110000000000,
31'b0000010000000000001000100000100,
31'b0000000000110000000010100000000,
31'b0000000000000000000101000010000,
31'b0110000000000000000000010101000,
31'b0100010000000000000100001000000,
31'b0100001000000010000000110000000,
31'b0100001000000000000000110000000,
31'b0000000100010000000001000000100,
31'b1000010000000000000001100010000,
31'b0000000001000000000010100000000,
31'b1000000000000000001100000000100,
31'b0010000000010000100010000001000,
31'b1100000000000100000000101000000,
31'b0010000000000001000000001000100,
31'b1100000000000000000000101000000,
31'b0000000100000000000001000000100,
31'b0000000100000010000001000000100,
31'b0000000100000100000001000000100,
31'b1000000100100000000000100100000,
31'b0010000000000000100010000001000,
31'b0010100000000000001000000000110,
31'b0010000000010001000000001000100,
31'b1100000000010000000000101000000,
31'b1000010000010000000110000000000,
31'b0101000010001000000000010000000,
31'b0000010000000000000000000110100,
31'b1000000100010000000000100100000,
31'b0101000010000010000000010000000,
31'b0101000010000000000000010000000,
31'b0010110000000000000010000000010,
31'b1100000000100000000000101000000,
31'b1000010000000000000110000000000,
31'b1000010000000010000110000000000,
31'b1000010000000100000110000000000,
31'b1000000100000000000000100100000,
31'b0010010010000000000000000000100,
31'b0101000010010000000000010000000,
31'b0010010010000100000000000000100,
31'b1101000000000000000100000000001,
31'b0000000010000000010000000000010,
31'b1001000000100000000000000100000,
31'b0001000000000000000001100000100,
31'b1001000000100100000000000100000,
31'b0001000000000000100000011000000,
31'b1001000000101000000000000100000,
31'b1000000010100000100000100000000,
31'b0110100000010000001000000000000,
31'b0001000101000000000010000000000,
31'b1001000000110000000000000100000,
31'b0100000100000000000001000000010,
31'b0110100000001000001000000000000,
31'b0001000101001000000010000000000,
31'b1101000100000000000000001000000,
31'b0110100000000010001000000000000,
31'b0110100000000000001000000000000,
31'b1001000000000010000000000100000,
31'b1001000000000000000000000100000,
31'b1001000000000110000000000100000,
31'b1001000000000100000000000100000,
31'b1001000000001010000000000100000,
31'b1001000000001000000000000100000,
31'b1000000010000000100000100000000,
31'b1001000000001100000000000100000,
31'b1010000011000000000000000001000,
31'b1001000000010000000000000100000,
31'b0100110000000000000000010000001,
31'b1001000000010100000000000100000,
31'b1001001001000000100000000000000,
31'b1000000000000000001000100001000,
31'b1010001000000000001000000100000,
31'b1011000010000000000000000010000,
31'b0001000100010000000010000000000,
31'b1010000000000001000010000000010,
31'b0100100010010000000000100000000,
31'b1010000000100000101000000000000,
31'b0001000100011000000010000000000,
31'b0010000000000101000000000010001,
31'b1000010000000000100000010000001,
31'b0010000000000001000000000010001,
31'b0001000100000000000010000000000,
31'b0001000100000010000010000000000,
31'b0100100010000000000000100000000,
31'b0100100010000010000000100000000,
31'b0001000100001000000010000000000,
31'b0101100000000000100000000100000,
31'b0100100010001000000000100000000,
31'b0100010100000000000000000000001,
31'b1010000010010000000000000001000,
31'b1001000001000000000000000100000,
31'b1010000000000010101000000000000,
31'b1010000000000000101000000000000,
31'b1001001000010000100000000000000,
31'b1010001000000000000000100010000,
31'b1000000000000000000000000111000,
31'b1010000000001000101000000000000,
31'b1010000010000000000000000001000,
31'b1010000010000010000000000001000,
31'b1010000010000100000000000001000,
31'b1010000000010000101000000000000,
31'b1001001000000000100000000000000,
31'b1001001000000010100000000000000,
31'b1001001000000100100000000000000,
31'b0100100000000000000001010000010,
31'b0000000000000000010000000000010,
31'b0000000000000010010000000000010,
31'b0000000000000100010000000000010,
31'b0000000000000110010000000000010,
31'b0000000000001000010000000000010,
31'b0000000000001010010000000000010,
31'b1000000000100000100000100000000,
31'b1001000000000000010001001000000,
31'b0000000000010000010000000000010,
31'b0000000001000001000000000100001,
31'b0100100001000000000000100000000,
31'b0100100001000010000000100000000,
31'b0000010001000000100100000000000,
31'b0000011000000000000000000000111,
31'b1010100000000000010100000000000,
31'b1011000000100000000000000010000,
31'b0000000000100000010000000000010,
31'b1001000010000000000000000100000,
31'b1000000000001000100000100000000,
31'b1001000010000100000000000100000,
31'b1000000000000100100000100000000,
31'b1001000010001000000000000100000,
31'b1000000000000000100000100000000,
31'b1000000000000010100000100000000,
31'b1010000001000000000000000001000,
31'b1010000001000010000000000001000,
31'b1010000001000100000000000001000,
31'b1011000000001000000000000010000,
31'b1010000001001000000000000001000,
31'b1011000000000100000000000010000,
31'b1000000000010000100000100000000,
31'b1011000000000000000000000010000,
31'b0000000001000000010000000000010,
31'b0000000001000010010000000000010,
31'b0100100000010000000000100000000,
31'b0100100000010010000000100000000,
31'b0000010000010000100100000000000,
31'b0000010000000000010001000000001,
31'b1100010000000000010000000001000,
31'b0011000000000000001001000000100,
31'b0000001000000000000001000000100,
31'b0000000000000001000000000100001,
31'b0100100000000000000000100000000,
31'b0100100000000010000000100000000,
31'b0000010000000000100100000000000,
31'b0000010000000010100100000000000,
31'b0100100000001000000000100000000,
31'b0100100000001010000000100000000,
31'b1010000000010000000000000001000,
31'b1010000000010010000000000001000,
31'b1010000000010100000000000001000,
31'b1010000010000000101000000000000,
31'b1010000000011000000000000001000,
31'b0100000100000001000000001000001,
31'b1000000001000000100000100000000,
31'b1001001000000000001000000001000,
31'b1010000000000000000000000001000,
31'b1010000000000010000000000001000,
31'b1010000000000100000000000001000,
31'b1000001000000000000000100100000,
31'b1010000000001000000000000001000,
31'b1010000000001010000000000001000,
31'b1010000000001100000000000001000,
31'b1011000001000000000000000010000,
31'b0001000001010000000010000000000,
31'b1001000100100000000000000100000,
31'b0100000000010000000001000000010,
31'b0100001000001001000100000000000,
31'b0001000100000000100000011000000,
31'b1101000000010000000000001000000,
31'b0100001000000011000100000000000,
31'b0100001000000001000100000000000,
31'b0001000001000000000010000000000,
31'b1000000000000000000000000001011,
31'b0100000000000000000001000000010,
31'b0100000000000010000001000000010,
31'b0001000001001000000010000000000,
31'b1101000000000000000000001000000,
31'b0100000000001000000001000000010,
31'b0000000000000000000010000011000,
31'b1001000100000010000000000100000,
31'b1001000100000000000000000100000,
31'b0100001000000000000000010011000,
31'b1001000100000100000000000100000,
31'b0010010000000000010001000000010,
31'b1100000000000000000100100000001,
31'b0000000010000001000000000010010,
31'b0100001000100001000100000000000,
31'b0010000000000001000000000100010,
31'b1001000100010000000000000100000,
31'b0100000000100000000001000000010,
31'b0100000010001000000000110000000,
31'b0010011001000000000000000000100,
31'b1101000000100000000000001000000,
31'b0100000010000010000000110000000,
31'b0100000010000000000000110000000,
31'b0001000000010000000010000000000,
31'b0010000000100000010000000000001,
31'b0100001000000000010000000000100,
31'b0100010000011000000000000000001,
31'b0001000000011000000010000000000,
31'b0101001000100000000000010000000,
31'b0100010000010010000000000000001,
31'b0100010000010000000000000000001,
31'b0001000000000000000010000000000,
31'b0001000000000010000010000000000,
31'b0001000000000100000010000000000,
31'b0100010000001000000000000000001,
31'b0001000000001000000010000000000,
31'b0100010000000100000000000000001,
31'b0100010000000010000000000000001,
31'b0100010000000000000000000000001,
31'b0010000000000010010000000000001,
31'b0010000000000000010000000000001,
31'b0110000000010000001000010000000,
31'b0010000000000100010000000000001,
31'b0101001000000010000000010000000,
31'b0101001000000000000000010000000,
31'b1000100000000000100001000000010,
31'b0101001000000100000000010000000,
31'b0001000000100000000010000000000,
31'b0010000000010000010000000000001,
31'b0110000000000000001000010000000,
31'b0110000000000010001000010000000,
31'b0010011000000000000000000000100,
31'b0101001000010000000000010000000,
31'b0110000000001000001000010000000,
31'b0100010000100000000000000000001,
31'b0000000100000000010000000000010,
31'b0010000000000000000010000101000,
31'b0000001000000000000010100000000,
31'b0000001000000010000010100000000,
31'b0000000100001000010000000000010,
31'b0010100000000000011001000000000,
31'b0000001000001000000010100000000,
31'b0100001010000001000100000000000,
31'b0001000011000000000010000000000,
31'b1011000000000001010000000000000,
31'b0100000010000000000001000000010,
31'b0100000010000010000001000000010,
31'b0001000011001000000010000000000,
31'b1101000010000000000000001000000,
31'b0100000010001000000001000000010,
31'b0100000000100000000000110000000,
31'b1000000000000001000010000000001,
31'b1001000110000000000000000100000,
31'b0000001000100000000010100000000,
31'b0100000000011000000000110000000,
31'b0000000000000101000000000010010,
31'b0100000001000001000000001000001,
31'b0000000000000001000000000010010,
31'b0100000000010000000000110000000,
31'b1010000101000000000000000001000,
31'b0100000000001100000000110000000,
31'b0100000010100000000001000000010,
31'b0100000000001000000000110000000,
31'b0100000000000110000000110000000,
31'b0100000000000100000000110000000,
31'b0100000000000010000000110000000,
31'b0100000000000000000000110000000,
31'b0001000010010000000010000000000,
31'b0010000010100000010000000000001,
31'b0001100000000000000000000000110,
31'b1000100000000000100000110000000,
31'b0001000010011000000010000000000,
31'b1100010000000000000100010000000,
31'b0011000000000000000010000110000,
31'b1100001000000000000000101000000,
31'b0001000010000000000010000000000,
31'b0001000010000010000010000000000,
31'b0100100100000000000000100000000,
31'b0100100100000010000000100000000,
31'b0001000010001000000010000000000,
31'b0101000000000001000100100000000,
31'b0100100100001000000000100000000,
31'b0100010010000000000000000000001,
31'b1010000100010000000000000001000,
31'b0010000010000000010000000000001,
31'b0001100000100000000000000000110,
31'b0010000010000100010000000000001,
31'b0100000000000011000000001000001,
31'b0100000000000001000000001000001,
31'b0000100000000000000000101100000,
31'b0100000001010000000000110000000,
31'b1010000100000000000000000001000,
31'b1010000100000010000000000001000,
31'b1010000100000100000000000001000,
31'b1010000000000000010100010000000,
31'b1010000100001000000000000001000,
31'b0100000001000100000000110000000,
31'b0100100000000000001000000000011,
31'b0100000001000000000000110000000,
31'b0101110000000000000000000000000,
31'b0000000010000000000100000100000,
31'b0101110000000100000000000000000,
31'b0000100000001000000010000000001,
31'b0101110000001000000000000000000,
31'b0000100000000100000010000000001,
31'b0001000000000000100100100000000,
31'b0000100000000000000010000000001,
31'b0101110000010000000000000000000,
31'b0010100000000000000000010000100,
31'b1000000000000010000000010100001,
31'b1000000000000000000000010100001,
31'b0010000101100000000000000000100,
31'b0010000000000100000100000010000,
31'b0010000000000010000100000010000,
31'b0010000000000000000100000010000,
31'b1001000000000000010100000000010,
31'b0000101000000000011000000000000,
31'b0010000000010001000000010001000,
31'b0000101000000100011000000000000,
31'b0010000101010000000000000000100,
31'b0000101000001000011000000000000,
31'b0010000000000000000011100000000,
31'b0000100000100000000010000000001,
31'b0010000101001000000000000000100,
31'b0010100000100000000000010000100,
31'b0010000000000001000000010001000,
31'b1000010000000000100000000011000,
31'b0010000101000000000000000000100,
31'b0100000110000000000100001000000,
31'b0000000000000000100000001000001,
31'b0010000000100000000100000010000,
31'b0110000000000000000000001100100,
31'b0000100000000000000001001001000,
31'b1100100000000000000000001000001,
31'b0000100001001000000010000000001,
31'b0010000100110000000000000000100,
31'b0000100001000100000010000000001,
31'b1001100000000000000000000001010,
31'b0000100001000000000010000000001,
31'b0011000000000000000100000001000,
31'b0011000000000010000100000001000,
31'b0011000000000100000100000001000,
31'b1100000000000000010000100010000,
31'b0010000100100000000000000000100,
31'b0100001100000100000000000000001,
31'b0100001100000010000000000000001,
31'b0100001100000000000000000000001,
31'b0010000100011000000000000000100,
31'b0000101001000000011000000000000,
31'b0000000100000000000010010000001,
31'b0000001000000000000000001100001,
31'b0010000100010000000000000000100,
31'b1010010000000000000000100010000,
31'b0010000100010100000000000000100,
31'b0000100010000000010000000101000,
31'b0010000100001000000000000000100,
31'b0100000100000000011010000000000,
31'b0010000100001100000000000000100,
31'b1100000000000000100010000000001,
31'b0010000100000000000000000000100,
31'b0100000000000000100000000010010,
31'b0010000100000100000000000000100,
31'b0100001100100000000000000000001,
31'b0000000000000010000100000100000,
31'b0000000000000000000100000100000,
31'b0000010100000000000010100000000,
31'b0000000000000100000100000100000,
31'b0000010000000001100000000000001,
31'b0000000000001000000100000100000,
31'b0001100100000001000000000100000,
31'b0000100010000000000010000000001,
31'b0000010001000000000001000000100,
31'b0000000000010000000100000100000,
31'b1000000100000000001001000100000,
31'b1000000000000000000010000010100,
31'b0000001001000000100100000000000,
31'b0000000000000000000000000000111,
31'b0110001000100000000000000000010,
31'b0010000010000000000100000010000,
31'b1000010000000000001000000010000,
31'b0000000000100000000100000100000,
31'b1000010000000100001000000010000,
31'b0000000001000000001011000000000,
31'b1000010000001000001000000010000,
31'b0000000000101000000100000100000,
31'b1100000000000000001001001000000,
31'b0000100010100000000010000000001,
31'b1000010000010000001000000010000,
31'b0000000100000000001000100000100,
31'b0110001000001000000000000000010,
31'b1000010001000000000000100100000,
31'b0110001000000100000000000000010,
31'b0100000100000000000100001000000,
31'b0110001000000000000000000000010,
31'b0110001000000010000000000000010,
31'b0000010000010000000001000000100,
31'b0000000001000000000100000100000,
31'b0000010101000000000010100000000,
31'b0000000001000100000100000100000,
31'b0000001000010000100100000000000,
31'b0000001000000000010001000000001,
31'b1100001000000000010000000001000,
31'b0000100011000000000010000000001,
31'b0000010000000000000001000000100,
31'b0000010000000010000001000000100,
31'b0000010000000100000001000000100,
31'b1000010000100000000000100100000,
31'b0000001000000000100100000000000,
31'b0000001000000010100100000000000,
31'b0100000000000000000000001010100,
31'b0100001110000000000000000000001,
31'b1000010001000000001000000010000,
31'b0000000001100000000100000100000,
31'b0000000100000000000000000110100,
31'b0000000000000000001011000000000,
31'b0010101000000000010000100000000,
31'b0000101000000000000110001000000,
31'b0110000000000000010001000000100,
31'b0000100000000000010000000101000,
31'b1000000100000000000110000000000,
31'b1000010000000100000000100100000,
31'b1000010000000010000000100100000,
31'b1000010000000000000000100100000,
31'b0010000110000000000000000000100,
31'b0100000101000000000100001000000,
31'b0110001001000000000000000000010,
31'b1001100000000001000010000000000,
31'b0101110100000000000000000000000,
31'b0000100000000001100000100000000,
31'b0100000000000000100000000100001,
31'b0100010000001001000100000000000,
31'b1010000000000000001001000010000,
31'b0101000010000000000000100000001,
31'b0100010000000011000100000000000,
31'b0100010000000001000100000000000,
31'b0011100000000001000000000010000,
31'b0010100100000000000000010000100,
31'b1000001000000000000010001000001,
31'b1001001000000000000001000010000,
31'b0010000001100000000000000000100,
31'b0100001001000100000000000000001,
31'b0100001001000010000000000000001,
31'b0100001001000000000000000000001,
31'b0010000001011000000000000000100,
31'b0010001000000000100000000100100,
31'b0000000001000000000010010000001,
31'b1001000000000000000000010001010,
31'b0010000001010000000000000000100,
31'b0101010001000000000000010000000,
31'b0010000100000000000011100000000,
31'b1100000000000000000000011000001,
31'b0010000001001000000000000000100,
31'b0010000000000001010100000000000,
31'b0010000100000001000000010001000,
31'b0011000000000000000000000011100,
31'b0010000001000000000000000000100,
31'b0100000010000000000100001000000,
31'b0010000001000100000000000000100,
31'b0100001001100000000000000000001,
31'b0111000000000000001000000000001,
31'b1000000010000000000001100010000,
31'b0100010000000000010000000000100,
31'b0100010000000010010000000000100,
31'b0010000000110000000000000000100,
31'b0101010000100000000000010000000,
31'b0100010000001000010000000000100,
31'b0100001000010000000000000000001,
31'b0010000000101000000000000000100,
31'b0100001000001100000000000000001,
31'b0100010000010000010000000000100,
31'b0100001000001000000000000000001,
31'b0010000000100000000000000000100,
31'b0100001000000100000000000000001,
31'b0100001000000010000000000000001,
31'b0100001000000000000000000000001,
31'b0010000000011000000000000000100,
31'b0101010000001000000000010000000,
31'b0000000000000000000010010000001,
31'b0001001000000000001000000000100,
31'b0010000000010000000000000000100,
31'b0101010000000000000000010000000,
31'b0010000000010100000000000000100,
31'b0101010000000100000000010000000,
31'b0010000000001000000000000000100,
31'b0100000000000000011010000000000,
31'b0010000000001100000000000000100,
31'b0100001000101000000000000000001,
31'b0010000000000000000000000000100,
31'b0010000000000010000000000000100,
31'b0010000000000100000000000000100,
31'b0100001000100000000000000000001,
31'b0000010000000100000010100000000,
31'b0000000100000000000100000100000,
31'b0000010000000000000010100000000,
31'b0000010000000010000010100000000,
31'b0101000000000010000000100000001,
31'b0101000000000000000000100000001,
31'b0001100000000001000000000100000,
31'b0101000000000100000000100000001,
31'b1000000001100000000110000000000,
31'b0000000100010000000100000100000,
31'b1000000000000000001001000100000,
31'b1000000100000000000010000010100,
31'b0110000000000000100000000010001,
31'b0100000000100000000100001000000,
31'b1000100000000000010010000001000,
31'b0100001011000000000000000000001,
31'b1000010100000000001000000010000,
31'b0000000100100000000100000100000,
31'b0000010000100000000010100000000,
31'b0000010000100010000010100000000,
31'b0111100000000000000001000000000,
31'b0100000000010000000100001000000,
31'b0011001000000000000000100000100,
31'b1101001000000001000000000000000,
31'b1000000001000000000110000000000,
31'b0000000000000000001000100000100,
31'b1000000001000100000110000000000,
31'b0000010000000000000101000010000,
31'b0100000000000010000100001000000,
31'b0100000000000000000100001000000,
31'b0110001100000000000000000000010,
31'b0100000000000100000100001000000,
31'b1000000000110000000110000000000,
31'b1000000000000000000001100010000,
31'b0000010001000000000010100000000,
31'b1000010000000000001100000000100,
31'b0010100000000001101000000000000,
31'b1100001000000000000100010000000,
31'b0010100000100000000010000000010,
31'b1100010000000000000000101000000,
31'b1000000000100000000110000000000,
31'b1000000000100010000110000000000,
31'b1000000001000000001001000100000,
31'b0100100000000000010000001001000,
31'b0010000010100000000000000000100,
31'b0100001010000100000000000000001,
31'b0100001010000010000000000000001,
31'b0100001010000000000000000000001,
31'b1000000000010000000110000000000,
31'b1000000000100000000001100010000,
31'b0000000000000000000000000110100,
31'b0000000100000000001011000000000,
31'b0010000010010000000000000000100,
31'b0101010010000000000000010000000,
31'b0010100000000000000010000000010,
31'b0010100000000010000010000000010,
31'b1000000000000000000110000000000,
31'b1000000000000010000110000000000,
31'b1000000000000100000110000000000,
31'b1000010100000000000000100100000,
31'b0010000010000000000000000000100,
31'b0100000001000000000100001000000,
31'b0010000010000100000000000000100,
31'b0100001010100000000000000000001,
31'b0001000000000000001100000010000,
31'b0000100000100000011000000000000,
31'b0010000010000000000100100001000,
31'b0000101000001000000010000000001,
31'b0001010000000000100000011000000,
31'b0000101000000100000010000000001,
31'b1000000001000000100000010000001,
31'b0000101000000000000010000000001,
31'b0001010101000000000010000000000,
31'b0010101000000000000000010000100,
31'b1000000100000000000010001000001,
31'b1001000100000000000001000010000,
31'b0000000100000000000000001010010,
31'b0110000000000000100000001000100,
31'b0110000010100000000000000000010,
31'b0100000101000000000000000000001,
31'b0100000000000000000000000110010,
31'b0000100000000000011000000000000,
31'b0100100000010000000000010000001,
31'b0000100000000100011000000000000,
31'b0110100000000000000010000000100,
31'b0000100000001000011000000000000,
31'b1100000000000000000010000100001,
31'b0000101000100000000010000000001,
31'b0100100000000100000000010000001,
31'b0000100000010000011000000000000,
31'b0100100000000000000000010000001,
31'b0100100000000010000000010000001,
31'b0110000010000100000000000000010,
31'b1001000000000001010001000000000,
31'b0110000010000000000000000000010,
31'b0110000010000010000000000000010,
31'b0001010100010000000010000000000,
31'b0000101000000000000001001001000,
31'b1010000000000001000000001001000,
31'b0000000000100000000000001100001,
31'b0000000100000000011000010000000,
31'b0000000010000000010001000000001,
31'b1000000000000000100000010000001,
31'b0000000000000000001100000001000,
31'b0001010100000000000010000000000,
31'b0100000100001100000000000000001,
31'b0100110010000000000000100000000,
31'b0100000100001000000000000000001,
31'b0000000010000000100100000000000,
31'b0100000100000100000000000000001,
31'b0100000100000010000000000000001,
31'b0100000100000000000000000000001,
31'b0100100000000001000000101000000,
31'b0000100001000000011000000000000,
31'b0000000000000010000000001100001,
31'b0000000000000000000000001100001,
31'b0010100010000000010000100000000,
31'b0000100010000000000110001000000,
31'b1000010000000000000000000111000,
31'b0000000000100000001100000001000,
31'b1010010010000000000000000001000,
31'b0100000000000100001000100000010,
31'b0100100001000000000000010000001,
31'b0100000000000000001000100000010,
31'b0010001100000000000000000000100,
31'b0100001000000000100000000010010,
31'b0110000011000000000000000000010,
31'b0100000100100000000000000000001,
31'b0000010000000000010000000000010,
31'b0000001000000000000100000100000,
31'b0010000000000000000100100001000,
31'b0000001000000100000100000100000,
31'b0000010000001000010000000000010,
31'b0000001000001000000100000100000,
31'b1100000001000000010000000001000,
31'b0000101010000000000010000000001,
31'b0000010000010000010000000000010,
31'b0000001000010000000100000100000,
31'b0110000000101000000000000000010,
31'b1001000000000001000000001100000,
31'b0000000001000000100100000000000,
31'b0000001000000000000000000000111,
31'b0110000000100000000000000000010,
31'b0110000000100010000000000000010,
31'b1100100000000000000100000000000,
31'b0000100010000000011000000000000,
31'b1100100000000100000100000000000,
31'b0000100010000100011000000000000,
31'b1100100000001000000100000000000,
31'b0000100010001000011000000000000,
31'b1000010000000000100000100000000,
31'b1101000100000001000000000000000,
31'b1100100000010000000100000000000,
31'b0000100100000000100100010000000,
31'b0110000000001000000000000000010,
31'b0110000000001010000000000000010,
31'b0110000000000100000000000000010,
31'b0110000000000110000000000000010,
31'b0110000000000000000000000000010,
31'b0110000000000010000000000000010,
31'b0000010001000000010000000000010,
31'b0000001001000000000100000100000,
31'b1100000000001000010000000001000,
31'b0000001001000100000100000100000,
31'b0000000000010000100100000000000,
31'b0000000000000000010001000000001,
31'b1100000000000000010000000001000,
31'b0000000010000000001100000001000,
31'b0000000000001000100100000000000,
31'b0000010000000001000000000100001,
31'b0100110000000000000000100000000,
31'b0100110000000010000000100000000,
31'b0000000000000000100100000000000,
31'b0000000000000010100100000000000,
31'b0000000000000100100100000000000,
31'b0100000110000000000000000000001,
31'b1100100001000000000100000000000,
31'b0000100011000000011000000000000,
31'b0001000100000001000010001000000,
31'b0000001000000000001011000000000,
31'b0010100000000000010000100000000,
31'b0000100000000000000110001000000,
31'b1100000000100000010000000001000,
31'b0000101000000000010000000101000,
31'b1010010000000000000000000001000,
31'b1010010000000010000000000001000,
31'b1010010000000100000000000001000,
31'b1010000000000000000010001000010,
31'b0000000000100000100100000000000,
31'b0010000000000000000000001010001,
31'b0110000001000000000000000000010,
31'b0110000001000010000000000000010,
31'b0001010001010000000010000000000,
31'b0010000010000000010000110000000,
31'b1010000000000000100001100000000,
31'b1001000000010000000001000010000,
31'b0000000001000000011000010000000,
31'b0100000001010100000000000000001,
31'b0100000001010010000000000000001,
31'b0100000001010000000000000000001,
31'b0001010001000000000010000000000,
31'b1001000000000100000001000010000,
31'b1000000000000000000010001000001,
31'b1001000000000000000001000010000,
31'b0000000000000000000000001010010,
31'b0100000001000100000000000000001,
31'b0100000001000010000000000000001,
31'b0100000001000000000000000000001,
31'b0100100000000000100001000001000,
31'b0010000000000000100000000100100,
31'b1001000000000000000110100000000,
31'b1000100000000000100000000000001,
31'b0010000000000000010001000000010,
31'b0010000000001000100000000100100,
31'b0011000010000000000000100000100,
31'b1101000010000001000000000000000,
31'b0010010000000001000000000100010,
31'b0010001000000001010100000000000,
31'b1000100000000000010101000000000,
31'b1001000000100000000001000010000,
31'b0010001001000000000000000000100,
31'b0100001010000000000100001000000,
31'b0110000110000000000000000000010,
31'b0100000001100000000000000000001,
31'b0001010000010000000010000000000,
31'b0110000000000000000010010000100,
31'b0100011000000000010000000000100,
31'b0100000000011000000000000000001,
31'b0000000000000000011000010000000,
31'b0100000000010100000000000000001,
31'b0100000000010010000000000000001,
31'b0100000000010000000000000000001,
31'b0001010000000000000010000000000,
31'b0100000000001100000000000000001,
31'b0100000000001010000000000000001,
31'b0100000000001000000000000000001,
31'b1000000000000000000001000001000,
31'b0100000000000100000000000000001,
31'b0100000000000010000000000000001,
31'b0100000000000000000000000000001,
31'b0010010000000010010000000000001,
31'b0010010000000000010000000000001,
31'b0001000000000010001000000000100,
31'b0001000000000000001000000000100,
31'b0010001000010000000000000000100,
31'b0101011000000000000000010000000,
31'b0111000000000000010010000000000,
31'b0100000000110000000000000000001,
31'b0010001000001000000000000000100,
31'b0100001000000000011010000000000,
31'b0110010000000000001000010000000,
31'b0100000000101000000000000000001,
31'b0010001000000000000000000000100,
31'b0100000000100100000000000000001,
31'b0100000000100010000000000000001,
31'b0100000000100000000000000000001,
31'b0000010100000000010000000000010,
31'b0010000000000000010000110000000,
31'b0010000000000000000000001100010,
31'b0010000000000100010000110000000,
31'b0000010100001000010000000000010,
31'b1100000001000000000100010000000,
31'b0011000000100000000000100000100,
31'b1101000000100001000000000000000,
31'b0001010011000000000010000000000,
31'b0010100000000001001000000100000,
31'b1000001000000000001001000100000,
31'b1001000010000000000001000010000,
31'b0000000101000000100100000000000,
31'b0100001000100000000100001000000,
31'b0110000100100000000000000000010,
31'b0100000011000000000000000000001,
31'b1100100100000000000100000000000,
31'b0010000010000000100000000100100,
31'b0011000000001000000000100000100,
31'b1101000000001001000000000000000,
31'b0011000000000100000000100000100,
31'b1101000000000101000000000000000,
31'b0011000000000000000000100000100,
31'b1101000000000001000000000000000,
31'b1000100000000000001000000001001,
31'b0000100000000000100100010000000,
31'b0110000100001000000000000000010,
31'b0100100000000000001001000000000,
31'b0110000100000100000000000000010,
31'b0100001000000000000100001000000,
31'b0110000100000000000000000000010,
31'b0000000000000000100000000010100,
31'b0001010010010000000010000000000,
31'b1100000000001000000100010000000,
31'b0010100000000001000000100010000,
31'b1100100000000000000000000010100,
31'b0000000100010000100100000000000,
31'b1100000000000000000100010000000,
31'b1100000100000000010000000001000,
31'b1000000000000000101001000000000,
31'b0001010010000000000010000000000,
31'b0100100000000000000110000100000,
31'b0100110100000000000000100000000,
31'b0100000010001000000000000000001,
31'b0000000100000000100100000000000,
31'b0100000010000100000000000000001,
31'b0100000010000010000000000000001,
31'b0100000010000000000000000000001,
31'b1100000000000001000000000011000,
31'b0010010010000000010000000000001,
31'b0001000000000001000010001000000,
31'b0001000010000000001000000000100,
31'b0010100100000000010000100000000,
31'b1100000000100000000100010000000,
31'b0011000001000000000000100000100,
31'b1101000001000001000000000000000,
31'b1000001000000000000110000000000,
31'b1000001000000010000110000000000,
31'b1000001000000100000110000000000,
31'b0100100001000000001001000000000,
31'b0010001010000000000000000000100,
31'b0100001001000000000100001000000,
31'b0110000101000000000000000000010,
31'b0100000010100000000000000000001,
31'b0110000000000000000000000000000,
31'b0110000000000010000000000000000,
31'b0110000000000100000000000000000,
31'b0110000000000110000000000000000,
31'b0110000000001000000000000000000,
31'b0110000000001010000000000000000,
31'b0110000000001100000000000000000,
31'b0110000000001110000000000000000,
31'b0110000000010000000000000000000,
31'b0110000000010010000000000000000,
31'b0110000000010100000000000000000,
31'b0110000000010110000000000000000,
31'b0110000000011000000000000000000,
31'b0110000000011010000000000000000,
31'b0000010000100000010000000000000,
31'b0101001000000000001000000000000,
31'b0110000000100000000000000000000,
31'b0110000000100010000000000000000,
31'b0000000000000001000001000100000,
31'b0000001000000000000000000000101,
31'b0110000000101000000000000000000,
31'b0110000000101010000000000000000,
31'b0000010000010000010000000000000,
31'b0000010000010010010000000000000,
31'b0110000000110000000000000000000,
31'b0110000000110010000000000000000,
31'b0000010000001000010000000000000,
31'b0000010000001010010000000000000,
31'b0000010000000100010000000000000,
31'b0010001000000000000010010000000,
31'b0000010000000000010000000000000,
31'b0000010000000010010000000000000,
31'b0110000001000000000000000000000,
31'b0110000001000010000000000000000,
31'b0110000001000100000000000000000,
31'b0110000001000110000000000000000,
31'b1000000000000000010100100000000,
31'b1010000000000000000010001000000,
31'b1010010000000000000000000001010,
31'b1010000000000100000010001000000,
31'b0110000001010000000000000000000,
31'b0110000001010010000000000000000,
31'b0110000001010100000000000000000,
31'b1000000100000001000011000000000,
31'b1010100000100000100000000000000,
31'b1010000000010000000010001000000,
31'b0100000000000000100000100001000,
31'b0101001001000000001000000000000,
31'b0110000001100000000000000000000,
31'b0110000001100010000000000000000,
31'b0000000000000000100100000000010,
31'b0000001001000000000000000000101,
31'b1010100000010000100000000000000,
31'b1010000000100000000010001000000,
31'b0000010001010000010000000000000,
31'b0000010001010010010000000000000,
31'b1100000000000000010000000001010,
31'b0001010000000000010000000011000,
31'b0000010001001000010000000000000,
31'b0000010000000001000100000000100,
31'b1010100000000000100000000000000,
31'b1010100000000010100000000000000,
31'b0000010001000000010000000000000,
31'b0000010001000010010000000000000,
31'b0110000010000000000000000000000,
31'b0110000010000010000000000000000,
31'b0110000010000100000000000000000,
31'b0110000010000110000000000000000,
31'b0000000000000001010000001000000,
31'b0100000001000000001000100000000,
31'b0100000000010000000000000110000,
31'b0100000001000100001000100000000,
31'b0110000010010000000000000000000,
31'b0110000010010010000000000000000,
31'b0100000000001000000000000110000,
31'b0110000000000000101000000001000,
31'b0100000000000100000000000110000,
31'b0100000001010000001000100000000,
31'b0100000000000000000000000110000,
31'b0100000000000010000000000110000,
31'b0110000010100000000000000000000,
31'b0110000010100010000000000000000,
31'b0000000100000000000000001010000,
31'b0000001010000000000000000000101,
31'b0100010100000000000001000000000,
31'b0100010100000010000001000000000,
31'b0000010010010000010000000000000,
31'b1000101000010000000000000010000,
31'b0110000010110000000000000000000,
31'b1000100000000000101000100000000,
31'b0000010010001000010000000000000,
31'b1000101000001000000000000010000,
31'b0010000000000001000001000010000,
31'b1000101000000100000000000010000,
31'b0000010010000000010000000000000,
31'b1000101000000000000000000010000,
31'b0110000011000000000000000000000,
31'b0000000000000000000100001000100,
31'b0110000011000100000000000000000,
31'b0100001000000000100000000010000,
31'b0100000000000010001000100000000,
31'b0100000000000000001000100000000,
31'b0100000001010000000000000110000,
31'b0100000000000100001000100000000,
31'b0110000011010000000000000000000,
31'b0101000000000000000000000101000,
31'b1001000000000000000001000100001,
31'b1001001000000001000000000000100,
31'b0100000001000100000000000110000,
31'b0100000000010000001000100000000,
31'b0100000001000000000000000110000,
31'b0100000001000010000000000110000,
31'b0110000011100000000000000000000,
31'b0100000100000000000000000000011,
31'b0000000101000000000000001010000,
31'b0100001000100000100000000010000,
31'b0100010101000000000001000000000,
31'b0100000000100000001000100000000,
31'b0001010100000000000010000000010,
31'b1100000100000000000010000010000,
31'b1001101000000000000000000001000,
31'b0001000000000000000000100000101,
31'b0000010011001000010000000000000,
31'b0011000000000001000001000001000,
31'b1010100010000000100000000000000,
31'b0100000100000000000100000100100,
31'b0000010011000000010000000000000,
31'b1010010000000001000010000000000,
31'b0110000100000000000000000000000,
31'b0110000100000010000000000000000,
31'b0110000100000100000000000000000,
31'b0110000100000110000000000000000,
31'b0110000100001000000000000000000,
31'b0110000100001010000000000000000,
31'b0110000100001100000000000000000,
31'b1000000001000000000000110001000,
31'b0000010000000001000000000010000,
31'b1010000000000000100000010000000,
31'b0010000010000000010001000000000,
31'b1010000000000100100000010000000,
31'b0010000000100000000000001100000,
31'b1010000000001000100000010000000,
31'b0100000000000001000001001000000,
31'b0101001100000000001000000000000,
31'b0110000100100000000000000000000,
31'b0110000100100010000000000000000,
31'b0000000010000000000000001010000,
31'b0000001100000000000000000000101,
31'b0100010010000000000001000000000,
31'b0110100001000000000000010000000,
31'b0000010100010000010000000000000,
31'b1000010010000000000000000001001,
31'b0010000000001000000000001100000,
31'b1010000000100000100000010000000,
31'b0000010100001000010000000000000,
31'b0000110000000000000000000011100,
31'b0010000000000000000000001100000,
31'b0010000000000010000000001100000,
31'b0000010100000000010000000000000,
31'b0000010100000010010000000000000,
31'b0110000101000000000000000000000,
31'b0110000101000010000000000000000,
31'b0110000101000100000000000000000,
31'b1000000000010001000011000000000,
31'b1010001000000000000000010100000,
31'b1010000100000000000010001000000,
31'b1000001000000000000110000000010,
31'b1000000000000000000000110001000,
31'b0010101000000000000010000000000,
31'b1010000001000000100000010000000,
31'b1000001010000000000000010010000,
31'b1000000000000001000011000000000,
31'b0010101000001000000010000000000,
31'b0001010000000101000000000001000,
31'b0100000100000000100000100001000,
31'b0001010000000001000000000001000,
31'b0110000101100000000000000000000,
31'b0100000010000000000000000000011,
31'b0000000100000000100100000000010,
31'b0110000000000000000100000010100,
31'b0110100000000010000000010000000,
31'b0110100000000000000000010000000,
31'b0001010010000000000010000000010,
31'b1100000010000000000010000010000,
31'b0010101000100000000010000000000,
31'b1110000000000000000010000100000,
31'b0001010000000000000100010010000,
31'b1100000000000000000100010000010,
31'b0010000001000000000000001100000,
31'b0110100000010000000000010000000,
31'b0001000000000000101000001000000,
31'b0001010000100001000000000001000,
31'b0110000110000000000000000000000,
31'b0110000110000010000000000000000,
31'b0000000000100000000000001010000,
31'b0010000000000000100100000000001,
31'b0100010000100000000001000000000,
31'b0100010000100010000001000000000,
31'b0010010000000001000000000100000,
31'b1000010000100000000000000001001,
31'b0010000000000100010001000000000,
31'b1010000010000000100000010000000,
31'b0010000000000000010001000000000,
31'b0010000000000010010001000000000,
31'b0100010000110000000001000000000,
31'b1001001000000000000000010001000,
31'b0100000100000000000000000110000,
31'b0100000100000010000000000110000,
31'b0000000000000100000000001010000,
31'b0100000001000000000000000000011,
31'b0000000000000000000000001010000,
31'b0000000000000010000000001010000,
31'b0100010000000000000001000000000,
31'b0100010000000010000001000000000,
31'b0000000000001000000000001010000,
31'b1000010000000000000000000001001,
31'b0100000000000001010000000100000,
31'b0100000001010000000000000000011,
31'b0000000000010000000000001010000,
31'b0000100000000000010000100000001,
31'b0100010000010000000001000000000,
31'b0100010000010010000001000000000,
31'b0000010110000000010000000000000,
31'b1000101100000000000000000010000,
31'b0110000111000000000000000000000,
31'b0100000000100000000000000000011,
31'b0010001000000000000000000000110,
31'b0100001100000000100000000010000,
31'b0100010001100000000001000000000,
31'b0100000100000000001000100000000,
31'b0010010001000001000000000100000,
31'b1100000000100000000010000010000,
31'b1000110000000000100001000000000,
31'b0101000100000000000000000101000,
31'b1000001000000000000000010010000,
31'b1000001000000010000000010010000,
31'b1000101000000000000100000000100,
31'b0001000000000000001000000000110,
31'b1100000000000000000101100000000,
31'b0010010000000000010000000000011,
31'b0100000000000010000000000000011,
31'b0100000000000000000000000000011,
31'b0000000001000000000000001010000,
31'b0100000000000100000000000000011,
31'b0100010001000000000001000000000,
31'b0001000000000000000000001001000,
31'b0001010000000000000010000000010,
31'b1100000000000000000010000010000,
31'b0100000001000001010000000100000,
31'b0100000000010000000000000000011,
31'b0000000001010000000000001010000,
31'b0100100000000000000000010110000,
31'b0100010001010000000001000000000,
31'b0100000000000000000100000100100,
31'b0001010000010000000010000000010,
31'b1100000000010000000010000010000,
31'b0110001000000000000000000000000,
31'b0110001000000010000000000000000,
31'b0110001000000100000000000000000,
31'b0000000000100000000000000000101,
31'b0110001000001000000000000000000,
31'b0110001000001010000000000000000,
31'b0110001000001100000000000000000,
31'b0101000000010000001000000000000,
31'b0110001000010000000000000000000,
31'b0110001000010010000000000000000,
31'b0110001000010100000000000000000,
31'b0101000000001000001000000000000,
31'b0110001000011000000000000000000,
31'b0101000000000100001000000000000,
31'b0101000000000010001000000000000,
31'b0101000000000000001000000000000,
31'b0110001000100000000000000000000,
31'b0000000000000100000000000000101,
31'b0000000000000010000000000000101,
31'b0000000000000000000000000000101,
31'b0110001000101000000000000000000,
31'b0010000000010000000010010000000,
31'b0000011000010000010000000000000,
31'b0000000000001000000000000000101,
31'b0110001000110000000000000000000,
31'b0010000000001000000010010000000,
31'b0000011000001000010000000000000,
31'b0000000000010000000000000000101,
31'b0010000000000010000010010000000,
31'b0010000000000000000010010000000,
31'b0000011000000000010000000000000,
31'b0000000000000000000100000100010,
31'b0110001001000000000000000000000,
31'b0110001001000010000000000000000,
31'b0110001001000100000000000000000,
31'b0100000010000000100000000010000,
31'b1010000100000000000000010100000,
31'b1010001000000000000010001000000,
31'b1000010000000000010000011000000,
31'b0101000001010000001000000000000,
31'b0100000000000000001000000011000,
31'b0110000000001000100000000100000,
31'b1001000000000000001010001000000,
31'b1001000010000001000000000000100,
31'b0110000000000010100000000100000,
31'b0110000000000000100000000100000,
31'b0101000001000010001000000000000,
31'b0101000001000000001000000000000,
31'b0110001001100000000000000000000,
31'b0010000100000000100000001000000,
31'b0000001000000000100100000000010,
31'b0000000001000000000000000000101,
31'b0001010010000000010000100000000,
31'b0010000100001000100000001000000,
31'b0000010000000000000001000000110,
31'b0000000001001000000000000000101,
31'b1110000000000000000000011000000,
31'b0010000100010000100000001000000,
31'b0000011001001000010000000000000,
31'b0000000001010000000000000000101,
31'b1010101000000000100000000000000,
31'b0010000001000000000010010000000,
31'b0000011001000000010000000000000,
31'b0000000000000001100001000000000,
31'b0110001010000000000000000000000,
31'b0110001010000010000000000000000,
31'b0110001010000100000000000000000,
31'b0100000001000000100000000010000,
31'b0101000000000000100000000001000,
31'b0101000000000010100000000001000,
31'b1001000000010000010100000000000,
31'b1001000000000000100001000000001,
31'b0110001010010000000000000000000,
31'b1000100100000001010000000000000,
31'b1001000000001000010100000000000,
31'b1001000001000001000000000000100,
31'b1001000000000100010100000000000,
31'b1001000100000000000000010001000,
31'b1001000000000000010100000000000,
31'b1000100000100000000000000010000,
31'b0110001010100000000000000000000,
31'b0010000000000000000100000010010,
31'b0000001100000000000000001010000,
31'b0000000010000000000000000000101,
31'b0101000000100000100000000001000,
31'b1000100000010100000000000010000,
31'b1000100000010010000000000010000,
31'b1000100000010000000000000010000,
31'b1001100001000000000000000001000,
31'b1000000000000000000100010000100,
31'b1000100000001010000000000010000,
31'b1000100000001000000000000010000,
31'b1000100000000110000000000010000,
31'b1000100000000100000000000010000,
31'b1000100000000010000000000010000,
31'b1000100000000000000000000010000,
31'b0110001011000000000000000000000,
31'b0100000000000100100000000010000,
31'b0100000000000010100000000010000,
31'b0100000000000000100000000010000,
31'b0101000001000000100000000001000,
31'b0100001000000000001000100000000,
31'b0110000000000000001000000101000,
31'b0100000000001000100000000010000,
31'b1001100000100000000000000001000,
31'b1001000000000101000000000000100,
31'b1000000100000000000000010010000,
31'b1001000000000001000000000000100,
31'b1000100100000000000100000000100,
31'b0110000010000000100000000100000,
31'b1001000001000000010100000000000,
31'b1001000000001001000000000000100,
31'b1001100000010000000000000001000,
31'b0100001100000000000000000000011,
31'b0110000000000000000100001000001,
31'b0100000000100000100000000010000,
31'b0001010000000000010000100000000,
31'b0100001000100000001000100000000,
31'b0011000000000000000100000001010,
31'b1100000000000001001000000000001,
31'b1001100000000000000000000001000,
31'b1001100000000010000000000001000,
31'b1001100000000100000000000001000,
31'b1001000000100001000000000000100,
31'b1000000000000001010000010000000,
31'b1000100001000100000000000010000,
31'b1000100001000010000000000010000,
31'b1000100001000000000000000010000,
31'b0110001100000000000000000000000,
31'b0110001100000010000000000000000,
31'b0110001100000100000000000000000,
31'b0100000000000000000100001000010,
31'b1101000000000000000101000000000,
31'b0001000010000000011001000000000,
31'b1001000000000000101000010000000,
31'b0001000000000000000100000001001,
31'b0010100001000000000010000000000,
31'b1010001000000000100000010000000,
31'b1000010000000000110010000000000,
31'b0101000100001000001000000000000,
31'b0010100001001000000010000000000,
31'b1110100000000000000000001000000,
31'b0101000100000010001000000000000,
31'b0101000100000000001000000000000,
31'b0110001100100000000000000000000,
31'b0010000001000000100000001000000,
31'b0000001010000000000000001010000,
31'b0000000100000000000000000000101,
31'b1110000000000000100010000000000,
31'b0010000100010000000010010000000,
31'b0000110010000000000000100000100,
31'b0000000100001000000000000000101,
31'b0010100001100000000010000000000,
31'b0010000100001000000010010000000,
31'b1000010000000000000000100010001,
31'b0000000100010000000000000000101,
31'b0010001000000000000000001100000,
31'b0010000100000000000010010000000,
31'b0000011100000000010000000000000,
31'b0000000000000000000000101001000,
31'b0000000000000000000100000010001,
31'b0010000000100000100000001000000,
31'b0010000010000000000000000000110,
31'b0100000110000000100000000010000,
31'b1010000000000000000000010100000,
31'b1010000000000010000000010100000,
31'b1000000000000000000110000000010,
31'b1000001000000000000000110001000,
31'b0010100000000000000010000000000,
31'b0010100000000010000010000000000,
31'b1000000010000000000000010010000,
31'b1000001000000001000011000000000,
31'b0010100000001000000010000000000,
31'b0110000100000000100000000100000,
31'b1000000010001000000000010010000,
31'b0101000101000000001000000000000,
31'b0010000000000010100000001000000,
31'b0010000000000000100000001000000,
31'b0010000010100000000000000000110,
31'b0010000000000100100000001000000,
31'b1010000000100000000000010100000,
31'b0010000000001000100000001000000,
31'b1100000000000001000001010000000,
31'b0010000000001100100000001000000,
31'b0010100000100000000010000000000,
31'b0010000000010000100000001000000,
31'b1100000000000000000010100001000,
31'b0010000000010100100000001000000,
31'b0010100000101000000010000000000,
31'b0010000101000000000010010000000,
31'b0101010000000000000001100000000,
31'b0000000100000001100001000000000,
31'b0110001110000000000000000000000,
31'b1000100000010001010000000000000,
31'b0010000001000000000000000000110,
31'b0100000101000000100000000010000,
31'b0101000100000000100000000001000,
31'b0001000000000000011001000000000,
31'b0010011000000001000000000100000,
31'b0010010000000000000001000000101,
31'b1000100000000011010000000000000,
31'b1000100000000001010000000000000,
31'b1000000001000000000000010010000,
31'b1000100000000101010000000000000,
31'b1001000000000010000000010001000,
31'b1001000000000000000000010001000,
31'b1001000100000000010100000000000,
31'b1001000000000100000000010001000,
31'b0100000000000000100100000000100,
31'b0100001001000000000000000000011,
31'b0000001000000000000000001010000,
31'b0000001000000010000000001010000,
31'b0100011000000000000001000000000,
31'b0100011000000010000001000000000,
31'b0000110000000000000000100000100,
31'b1000100100010000000000000010000,
31'b1001000000000001000100000010000,
31'b1000100000100001010000000000000,
31'b1000000000000000010000000001100,
31'b1000100100001000000000000010000,
31'b0100011000010000000001000000000,
31'b1001000000100000000000010001000,
31'b1000100100000010000000000010000,
31'b1000100100000000000000000010000,
31'b0010000000000100000000000000110,
31'b0100001000100000000000000000011,
31'b0010000000000000000000000000110,
31'b0100000100000000100000000010000,
31'b1010000010000000000000010100000,
31'b0100001100000000001000100000000,
31'b0010000000001000000000000000110,
31'b0100000100001000100000000010000,
31'b1000000000000100000000010010000,
31'b1000100001000001010000000000000,
31'b1000000000000000000000010010000,
31'b1000000000000010000000010010000,
31'b1000100000000000000100000000100,
31'b1001000001000000000000010001000,
31'b1000000000001000000000010010000,
31'b1000000000100001000100000001000,
31'b0100001000000010000000000000011,
31'b0100001000000000000000000000011,
31'b0010000000100000000000000000110,
31'b0100001000000100000000000000011,
31'b0100011001000000000001000000000,
31'b0100000000000001110000000000000,
31'b0011000000000000000000101100000,
31'b1100001000000000000010000010000,
31'b1001100100000000000000000001000,
31'b0100010000000000100001000100000,
31'b1000000000100000000000010010000,
31'b1000000000100010000000010010000,
31'b1000100000100000000100000000100,
31'b1001000000000000010000000010100,
31'b1000000000101000000000010010000,
31'b1000000000000001000100000001000,
31'b0110010000000000000000000000000,
31'b0110010000000010000000000000000,
31'b0110010000000100000000000000000,
31'b0110010000000110000000000000000,
31'b0110010000001000000000000000000,
31'b0110010000001010000000000000000,
31'b0000000000110000010000000000000,
31'b0011000000000000000010000000001,
31'b0000000100000001000000000010000,
31'b0001000000000000000000010000100,
31'b0000000000101000010000000000000,
31'b0001000000000100000000010000100,
31'b0000000000100100010000000000000,
31'b0001000000001000000000010000100,
31'b0000000000100000010000000000000,
31'b0000000000100010010000000000000,
31'b0110010000100000000000000000000,
31'b0110010000100010000000000000000,
31'b0000000000011000010000000000000,
31'b0000011000000000000000000000101,
31'b0000000000010100010000000000000,
31'b0100000000000000001000010000001,
31'b0000000000010000010000000000000,
31'b0000000000010010010000000000000,
31'b0000000000001100010000000000000,
31'b0001000000100000000000010000100,
31'b0000000000001000010000000000000,
31'b0000000000001010010000000000000,
31'b0000000000000100010000000000000,
31'b0000000000000110010000000000000,
31'b0000000000000000010000000000000,
31'b0000000000000010010000000000000,
31'b0110010001000000000000000000000,
31'b0110010001000010000000000000000,
31'b1100100000000000110000000000000,
31'b0000100100010000010000010000000,
31'b1010000000000100000000000001010,
31'b1010010000000000000010001000000,
31'b1010000000000000000000000001010,
31'b1010000000000010000000000001010,
31'b0000100000000000000100000001000,
31'b0001000001000000000000010000100,
31'b0000100000000100000100000001000,
31'b0000100100000000010000010000000,
31'b0000100000001000000100000001000,
31'b0001000100000101000000000001000,
31'b0000000001100000010000000000000,
31'b0001000100000001000000000001000,
31'b0110010001100000000000000000000,
31'b1001001000000000000000001000100,
31'b0000010000000000100100000000010,
31'b0000001000000000110000000100000,
31'b0100100000000000000000100000010,
31'b0100100000000010000000100000010,
31'b0000000001010000010000000000000,
31'b0000000001010010010000000000000,
31'b0000100000100000000100000001000,
31'b0001000000000000010000000011000,
31'b0000000001001000010000000000000,
31'b0000000000000001000100000000100,
31'b0000000001000100010000000000000,
31'b0000100000000001000000010010000,
31'b0000000001000000010000000000000,
31'b0000000001000010010000000000000,
31'b0110010010000000000000000000000,
31'b0110010010000010000000000000000,
31'b0110010010000100000000000000000,
31'b1001000000000000000100000000101,
31'b0100000100100000000001000000000,
31'b0100010001000000001000100000000,
31'b0010000100000001000000000100000,
31'b1001000000010000000000000100010,
31'b0000000000000000000001001100000,
31'b0001000010000000000000010000100,
31'b0000000010101000010000000000000,
31'b1001000000001000000000000100010,
31'b0000000010100100010000000000000,
31'b1001000000000100000000000100010,
31'b0000000010100000010000000000000,
31'b1001000000000000000000000100010,
31'b0100000100001000000001000000000,
31'b0110100000000000001000000000010,
31'b0000010100000000000000001010000,
31'b1000000100001000000000000001001,
31'b0100000100000000000001000000000,
31'b0100000100000010000001000000000,
31'b0000000010010000010000000000000,
31'b1000000100000000000000000001001,
31'b0000000010001100010000000000000,
31'b1000000000001000100001010000000,
31'b0000000010001000010000000000000,
31'b1000000000000000000000101000100,
31'b0000000010000100010000000000000,
31'b1000000000000000100001010000000,
31'b0000000010000000010000000000000,
31'b0000000010000010010000000000000,
31'b0110010011000000000000000000000,
31'b0100100000000000000001010000000,
31'b1001001000000000100000000000010,
31'b0000100000000000101100000000000,
31'b0100010000000010001000100000000,
31'b0100010000000000001000100000000,
31'b1010000010000000000000000001010,
31'b0100010000000100001000100000000,
31'b0000100010000000000100000001000,
31'b0101010000000000000000000101000,
31'b0000100010000100000100000001000,
31'b0010001100000001100000000000000,
31'b0000101000100000000011000000000,
31'b1100000000000000000011000100000,
31'b0000000011100000010000000000000,
31'b1010000000100001000010000000000,
31'b1001000100000000000000000010001,
31'b1000000100000000000011001000000,
31'b0001000100001000000010000000010,
31'b0010100000000001000000010100000,
31'b0100000101000000000001000000000,
31'b0100010000100000001000100000000,
31'b0001000100000000000010000000010,
31'b1010000000010001000010000000000,
31'b0000101000001000000011000000000,
31'b0010000000000100011000100000000,
31'b0000000011001000010000000000000,
31'b0010000000000000011000100000000,
31'b0000101000000000000011000000000,
31'b1010000000000101000010000000000,
31'b0000000011000000010000000000000,
31'b1010000000000001000010000000000,
31'b0000000000010001000000000010000,
31'b0100000000000000000000110000010,
31'b0100000000000000010000001100000,
31'b0100000000000100000000110000010,
31'b0100000010100000000001000000000,
31'b0100000010100010000001000000000,
31'b0010000010000001000000000100000,
31'b1000000010100000000000000001001,
31'b0000000000000001000000000010000,
31'b0000000000000011000000000010000,
31'b0000000000000101000000000010000,
31'b0000100001000000010000010000000,
31'b0000000000001001000000000010000,
31'b0000000000100000000100010001000,
31'b0000000100100000010000000000000,
31'b0001000001000001000000000001000,
31'b0100000010001000000001000000000,
31'b0100000010001010000001000000000,
31'b0000010010000000000000001010000,
31'b1000101000000000010000001000000,
31'b0100000010000000000001000000000,
31'b0100000010000010000001000000000,
31'b0000000100010000010000000000000,
31'b1000000010000000000000000001001,
31'b0000000000100001000000000010000,
31'b0000000000100011000000000010000,
31'b0000000100001000010000000000000,
31'b0000100000000000000000000011100,
31'b0000000100000100010000000000000,
31'b0000000000000000000100010001000,
31'b0000000100000000010000000000000,
31'b0000000100000010010000000000000,
31'b0100100000000000001000000000001,
31'b0100100000000010001000000000001,
31'b0100100000000100001000000000001,
31'b0000100000010000010000010000000,
31'b0100100000001000001000000000001,
31'b1000001000000000000100001001000,
31'b1010000100000000000000000001010,
31'b1000000000000000010010000100000,
31'b0000000001000001000000000010000,
31'b0000100000000100010000010000000,
31'b0000100000000010010000010000000,
31'b0000100000000000010000010000000,
31'b0001100000100000000000000000100,
31'b0001000000000101000000000001000,
31'b0001000000000011000000000001000,
31'b0001000000000001000000000001000,
31'b1001000010000000000000000010001,
31'b1000001000000000001000000100001,
31'b0001000010001000000010000000010,
31'b0010101000000000001000000000100,
31'b0100000011000000000001000000000,
31'b0110110000000000000000010000000,
31'b0001000010000000000010000000010,
31'b1000000011000000000000000001001,
31'b0001100000001000000000000000100,
31'b0001100000001010000000000000100,
31'b0001000000000000000100010010000,
31'b0000100000100000010000010000000,
31'b0001100000000000000000000000100,
31'b0001100000000010000000000000100,
31'b0000000101000000010000000000000,
31'b0001000000100001000000000001000,
31'b0100000000101000000001000000000,
31'b0100000010000000000000110000010,
31'b0010000000001001000000000100000,
31'b1000000000101000000000000001001,
31'b0100000000100000000001000000000,
31'b0100000000100010000001000000000,
31'b0010000000000001000000000100000,
31'b1000000000100000000000000001001,
31'b0000000010000001000000000010000,
31'b0000001000000000000011010000000,
31'b0010010000000000010001000000000,
31'b0010010000000010010001000000000,
31'b0100000000110000000001000000000,
31'b0100000000110010000001000000000,
31'b0010000000010001000000000100000,
31'b1001000100000000000000000100010,
31'b0100000000001000000001000000000,
31'b0100000000001010000001000000000,
31'b0000010000000000000000001010000,
31'b1000000000001000000000000001001,
31'b0100000000000000000001000000000,
31'b0100000000000010000001000000000,
31'b0100000000000100000001000000000,
31'b1000000000000000000000000001001,
31'b0100000000011000000001000000000,
31'b0100001000000001000100000000010,
31'b0000010000010000000000001010000,
31'b1000000100000000000000101000100,
31'b0100000000010000000001000000000,
31'b0100000000010010000001000000000,
31'b0000000110000000010000000000000,
31'b1000000000010000000000000001001,
31'b1001000000100000000000000010001,
31'b1000100000000000010100000000001,
31'b0010011000000000000000000000110,
31'b0010001000010001100000000000000,
31'b0100000001100000000001000000000,
31'b0100010100000000001000100000000,
31'b0010000001000001000000000100000,
31'b1000000010000000010010000100000,
31'b1000100000000000100001000000000,
31'b1010000000000000010010000010000,
31'b1000100000000100100001000000000,
31'b0010001000000001100000000000000,
31'b1100000000000000001000000010100,
31'b0010000000000100010000000000011,
31'b0010000001010001000000000100000,
31'b0010000000000000010000000000011,
31'b1001000000000000000000000010001,
31'b1000000000000000000011001000000,
31'b0001000000001000000010000000010,
31'b1000000001001000000000000001001,
31'b0100000001000000000001000000000,
31'b0100000001000010000001000000000,
31'b0001000000000000000010000000010,
31'b1000000001000000000000000001001,
31'b1001000000010000000000000010001,
31'b1010000000000000100000100000001,
31'b0001000010000000000100010010000,
31'b0010001000100001100000000000000,
31'b0100000001010000000001000000000,
31'b0100010000000000000100000100100,
31'b0001000000010000000010000000010,
31'b1010000100000001000010000000000,
31'b0110011000000000000000000000000,
31'b0110011000000010000000000000000,
31'b0110011000000100000000000000000,
31'b0100000000000000010010010000000,
31'b0110011000001000000000000000000,
31'b1000100000000001000000001010000,
31'b0010000000000000001000010000100,
31'b0101010000010000001000000000000,
31'b0000000000000000001010000000001,
31'b0001001000000000000000010000100,
31'b0000001000101000010000000000000,
31'b0101010000001000001000000000000,
31'b0000001000100100010000000000000,
31'b0110000000000000010000000000101,
31'b0000001000100000010000000000000,
31'b0101010000000000001000000000000,
31'b0110011000100000000000000000000,
31'b0011000000000000011000000000000,
31'b0000010000000010000000000000101,
31'b0000010000000000000000000000101,
31'b0101000000000000000010000000100,
31'b0101000000000010000010000000100,
31'b0000001000010000010000000000000,
31'b0000010000001000000000000000101,
31'b0000001000001100010000000000000,
31'b0011000000010000011000000000000,
31'b0000001000001000010000000000000,
31'b0000010000010000000000000000101,
31'b0000001000000100010000000000000,
31'b0010010000000000000010010000000,
31'b0000001000000000010000000000000,
31'b0000001000000010010000000000000,
31'b0110011001000000000000000000000,
31'b1001000000100000000000001000100,
31'b1001000010000000100000000000010,
31'b0000000010000000000000110000100,
31'b1000000000000100010000011000000,
31'b1000000000000000000000100100010,
31'b1000000000000000010000011000000,
31'b1000000000000100000000100100010,
31'b0000101000000000000100000001000,
31'b1001000000000000001000000001010,
31'b0000101000000100000100000001000,
31'b0010100000000000000100100100000,
31'b0000101000001000000100000001000,
31'b1100000000000000001000001000001,
31'b0000001001100000010000000000000,
31'b0101010001000000001000000000000,
31'b1001000000000010000000001000100,
31'b1001000000000000000000001000100,
31'b0000000000001000000001000000110,
31'b0000000000000000110000000100000,
31'b0001000010000000010000100000000,
31'b1001000000001000000000001000100,
31'b0000000000000000000001000000110,
31'b0000000000001000110000000100000,
31'b0000101000100000000100000001000,
31'b1100000000000000000100000101000,
31'b0000001001001000010000000000000,
31'b0000001000000001000100000000100,
31'b0000100010000000000011000000000,
31'b0010010001000000000010010000000,
31'b0000001001000000010000000000000,
31'b0000010000000001100001000000000,
31'b1100000000000000100011000000000,
31'b0000000100010000000011010000000,
31'b1001000001000000100000000000010,
31'b0000000001000000000000110000100,
31'b0101010000000000100000000001000,
31'b0000000100000001000000100001000,
31'b0010001100000001000000000100000,
31'b0010000100000000000001000000101,
31'b0000001000000000000001001100000,
31'b0000000100000000000011010000000,
31'b0000100000100000000000001001001,
31'b0010000101000001100000000000000,
31'b0000100001100000000011000000000,
31'b0010000001000000000010100000001,
31'b0000100000000000001100000100000,
31'b1001001000000000000000000100010,
31'b1111000000000000000100000000000,
31'b0011000010000000011000000000000,
31'b0000100100001000000000100000100,
31'b0000010010000000000000000000101,
31'b0100001100000000000001000000000,
31'b0101000000000001001000001000000,
31'b0000100100000000000000100000100,
31'b1000110000010000000000000010000,
31'b0000100001001000000011000000000,
31'b1100100000000000000001001000000,
31'b0000100000000000000000001001001,
31'b1000110000001000000000000010000,
31'b0000100001000000000011000000000,
31'b1000110000000100000000000010000,
31'b0000001010000000010000000000000,
31'b1000110000000000000000000010000,
31'b1001000000000100100000000000010,
31'b0000000000001000100001001000000,
31'b1001000000000000100000000000010,
31'b0000000000000000000000110000100,
31'b0001000000100000010000100000000,
31'b0000000000000000100001001000000,
31'b1001000000001000100000000000010,
31'b0000000000001000000000110000100,
31'b0000101010000000000100000001000,
31'b0010000100000101100000000000000,
31'b1001000000010000100000000000010,
31'b0010000100000001100000000000000,
31'b0000100000100000000011000000000,
31'b0010000000000000000010100000001,
31'b0000100001000000001100000100000,
31'b0010000100001001100000000000000,
31'b1000000000000000000001010100000,
31'b1001000010000000000000001000100,
31'b1001000000100000100000000000010,
31'b0000000010000000110000000100000,
31'b0001000000000000010000100000000,
31'b0001000000000010010000100000000,
31'b0001000000000100010000100000000,
31'b0001000000000110010000100000000,
31'b0000100000001000000011000000000,
31'b0100100000000000000000000011010,
31'b0000100001000000000000001001001,
31'b0010001000000000011000100000000,
31'b0000100000000000000011000000000,
31'b0010000000000000110000000010000,
31'b0000100000000100000011000000000,
31'b1010001000000001000010000000000,
31'b0100000000000000000110000001000,
31'b0100001000000000000000110000010,
31'b1001000000000000000100001010000,
31'b1000100000100000010000001000000,
31'b0100001010100000000001000000000,
31'b0000000010000001000000100001000,
31'b0010001010000001000000000100000,
31'b0011000000000001001000000010000,
31'b0000001000000001000000000010000,
31'b0000001000000011000000000010000,
31'b1000000000000000110010000000000,
31'b1010100000000000000001000010000,
31'b0000001000001001000000000010000,
31'b0000001000100000000100010001000,
31'b0000001100100000010000000000000,
31'b0101010100000000001000000000000,
31'b0100001010001000000001000000000,
31'b1000100000000100010000001000000,
31'b1000100000000010010000001000000,
31'b1000100000000000010000001000000,
31'b0100001010000000000001000000000,
31'b0100001010000010000001000000000,
31'b0000100010000000000000100000100,
31'b1000100000001000010000001000000,
31'b0000001000100001000000000010000,
31'b0100000010000001000100000000010,
31'b1000000000000000000000100010001,
31'b1000100000010000010000001000000,
31'b0000000000000000000010100000010,
31'b0000001000000000000100010001000,
31'b0000001100000000010000000000000,
31'b0000010000000000000000101001000,
31'b0010000000000001001000000001000,
31'b1000000000100000001000000100001,
31'b0010010010000000000000000000110,
31'b0010100000100000001000000000100,
31'b1010010000000000000000010100000,
31'b1000000000000000000100001001000,
31'b1000010000000000000110000000010,
31'b1000001000000000010010000100000,
31'b0010110000000000000010000000000,
31'b0010110000000010000010000000000,
31'b1000010010000000000000010010000,
31'b0010000010000001100000000000000,
31'b0011000000000001000000100100000,
31'b1101000000000000000000000100100,
31'b0101000000100000000001100000000,
31'b0100000000000000110000001000000,
31'b1000000000000010001000000100001,
31'b1000000000000000001000000100001,
31'b0100100000001000010010000000000,
31'b0010100000000000001000000000100,
31'b0100100000000100010010000000000,
31'b1000000000100000000100001001000,
31'b0100100000000000010010000000000,
31'b0110000000000000100001000010000,
31'b0010110000100000000010000000000,
31'b1100000000000000000000101000010,
31'b1100000000000000010000010100000,
31'b0010100000010000001000000000100,
31'b0001101000000000000000000000100,
31'b1001000000000000000000100001001,
31'b0101000000000000000001100000000,
31'b0101000000000010000001100000000,
31'b0100001000101000000001000000000,
31'b0000000000010000000011010000000,
31'b0010010001000000000000000000110,
31'b0010000001010001100000000000000,
31'b0100001000100000000001000000000,
31'b0000000000000001000000100001000,
31'b0010001000000001000000000100000,
31'b0010000000000000000001000000101,
31'b0000001010000001000000000010000,
31'b0000000000000000000011010000000,
31'b1000010001000000000000010010000,
31'b0010000001000001100000000000000,
31'b0100001000110000000001000000000,
31'b0000000000010001000000100001000,
31'b0010001000010001000000000100000,
31'b0010000001001001100000000000000,
31'b0100001000001000000001000000000,
31'b0100001000001010000001000000000,
31'b0000100000001000000000100000100,
31'b1000100010000000010000001000000,
31'b0100001000000000000001000000000,
31'b0100001000000010000001000000000,
31'b0000100000000000000000100000100,
31'b1000001000000000000000000001001,
31'b0100001000011000000001000000000,
31'b0100000000000001000100000000010,
31'b1000010000000000010000000001100,
31'b0111000000000000001001000000000,
31'b0100001000010000000001000000000,
31'b0100001000010010000001000000000,
31'b0000100000010000000000100000100,
31'b1000110100000000000000000010000,
31'b0010010000000100000000000000110,
31'b0010000000010101100000000000000,
31'b0010010000000000000000000000110,
31'b0010000000010001100000000000000,
31'b0100001001100000000001000000000,
31'b0000000100000000100001001000000,
31'b0010010000001000000000000000110,
31'b0010000001000000000001000000101,
31'b1000101000000000100001000000000,
31'b0010000000000101100000000000000,
31'b1000010000000000000000010010000,
31'b0010000000000001100000000000000,
31'b1100000000000000000001011000000,
31'b0010000100000000000010100000001,
31'b1000010000001000000000010010000,
31'b0010000000001001100000000000000,
31'b1001001000000000000000000010001,
31'b1000001000000000000011001000000,
31'b0010100000000001000010001000000,
31'b0010100010000000001000000000100,
31'b0100001001000000000001000000000,
31'b0100010000000001110000000000000,
31'b0001001000000000000010000000010,
31'b1000100000000000001110000000000,
31'b0100000000001000010000000000110,
31'b0100000000000000100001000100000,
31'b1000010000100000000000010010000,
31'b0010000000100001100000000000000,
31'b0100000000000000010000000000110,
31'b0100000000001000100001000100000,
31'b0101000010000000000001100000000,
31'b1010000000000000001000000010001,
31'b0110100000000000000000000000000,
31'b0110100000000010000000000000000,
31'b1000000000100000000000100001000,
31'b1100001000000001000001000000000,
31'b0110100000001000000000000000000,
31'b0110100000001010000000000000000,
31'b1100000000010000000100000000010,
31'b0001010000010000000100000010000,
31'b0110100000010000000000000000000,
31'b0110100000010010000000000000000,
31'b1100000000001000000100000000010,
31'b0001010000001000000100000010000,
31'b1100000000000100000100000000010,
31'b0001010000000100000100000010000,
31'b1100000000000000000100000000010,
31'b0001010000000000000100000010000,
31'b1000000000000100000000100001000,
31'b1010001000000000000000000100000,
31'b1000000000000000000000100001000,
31'b1000000000000010000000100001000,
31'b1010000001010000100000000000000,
31'b1010001000001000000000000100000,
31'b1000000000001000000000100001000,
31'b1000001010010000000000000010000,
31'b1010000001001000100000000000000,
31'b1010001000010000000000000100000,
31'b1000000000010000000000100001000,
31'b1000001010001000000000000010000,
31'b1010000001000000100000000000000,
31'b1010000001000010100000000000000,
31'b0000110000000000010000000000000,
31'b1000001010000000000000000010000,
31'b0110100001000000000000000000000,
31'b0110100001000010000000000000000,
31'b1100010000000000110000000000000,
31'b0001000100001000001010000000000,
31'b1010000000110000100000000000000,
31'b1010100000000000000010001000000,
31'b0001000100000010001010000000000,
31'b0001000100000000001010000000000,
31'b0000010000000000000100000001000,
31'b0010000000000000000000011100000,
31'b0010000000000000010000100000010,
31'b0000010100000000010000010000000,
31'b1010000000100000100000000000000,
31'b1010000000100010100000000000000,
31'b1100000001000000000100000000010,
31'b0001010001000000000100000010000,
31'b1010000000011000100000000000000,
31'b1010001001000000000000000100000,
31'b1000000001000000000000100001000,
31'b1001001000000000101000000000000,
31'b1010000000010000100000000000000,
31'b1001000000000000000000100010000,
31'b1010000000010100100000000000000,
31'b1010000010000000001000000001000,
31'b1010000000001000100000000000000,
31'b1010000000001010100000000000000,
31'b1010000000001100100000000000000,
31'b0100000100000000000010000000101,
31'b1010000000000000100000000000000,
31'b1010000000000010100000000000000,
31'b1010000000000100100000000000000,
31'b1010000000000110100000000000000,
31'b0110100010000000000000000000000,
31'b0110100010000010000000000000000,
31'b1100000000000000000010010010000,
31'b0001010000000000000010010000010,
31'b0100000000000000000000010000011,
31'b0100100001000000001000100000000,
31'b0100100000010000000000000110000,
31'b0000000001000000000000011010000,
31'b0110100010010000000000000000000,
31'b1000001100000001010000000000000,
31'b0110000000000000000010000000110,
31'b0000000100000000100010000010000,
31'b0100100000000100000000000110000,
31'b0000000000000100011000000000010,
31'b0100100000000000000000000110000,
31'b0000000000000000011000000000010,
31'b1011000000000000001000000010000,
31'b1010001010000000000000000100000,
31'b1000000010000000000000100001000,
31'b1000001000011000000000000010000,
31'b0100110100000000000001000000000,
31'b1001000000000000100000000101000,
31'b1000001000010010000000000010000,
31'b1000001000010000000000000010000,
31'b1001001001000000000000000001000,
31'b1000000000000000101000100000000,
31'b1000001000001010000000000010000,
31'b1000001000001000000000000010000,
31'b1010000011000000100000000000000,
31'b1000001000000100000000000010000,
31'b1000001000000010000000000010000,
31'b1000001000000000000000000010000,
31'b0110100011000000000000000000000,
31'b0100010000000000000001010000000,
31'b1000010000000000000000010001001,
31'b0000010000000000101100000000000,
31'b0100100000000010001000100000000,
31'b0100100000000000001000100000000,
31'b0000000000000010000000011010000,
31'b0000000000000000000000011010000,
31'b0011000000000000000001000000100,
31'b0101100000000000000000000101000,
31'b0011000000000100000001000000100,
31'b0000010110000000010000010000000,
31'b1010000010100000100000000000000,
31'b0100100000010000001000100000000,
31'b0100100001000000000000000110000,
31'b0000000001000000011000000000010,
31'b1001001000010000000000000001000,
31'b0100100100000000000000000000011,
31'b1000000000000000100000000110000,
31'b1010000000001000001000000001000,
31'b1010000010010000100000000000000,
31'b1010000000000100001000000001000,
31'b1010000000000010001000000001000,
31'b1010000000000000001000000001000,
31'b1001001000000000000000000001000,
31'b1001001000000010000000000001000,
31'b1001001000000100000000000001000,
31'b1011000000000000000000100100000,
31'b1010000010000000100000000000000,
31'b1010000010000010100000000000000,
31'b1010000010000100100000000000000,
31'b1000001001000000000000000010000,
31'b0110100100000000000000000000000,
31'b0110100100000010000000000000000,
31'b1101000000000000001000001000000,
31'b0001000010000000010100001000000,
31'b0110100100001000000000000000000,
31'b0100000000000000001001000000010,
31'b1001000000000000000100100000100,
31'b0001000001000000001010000000000,
31'b0010001001000000000010000000000,
31'b1010100000000000100000010000000,
31'b0010100010000000010001000000000,
31'b0000010001000000010000010000000,
31'b0010100000100000000000001100000,
31'b1110001000000000000000001000000,
31'b1100000100000000000100000000010,
31'b0001010100000000000100000010000,
31'b1010000000000000000010011000000,
31'b1010001100000000000000000100000,
31'b1000000100000000000000100001000,
31'b1000011000000000010000001000000,
31'b0110000001000010000000010000000,
31'b0110000001000000000000010000000,
31'b1000000100001000000000100001000,
31'b0110000001000100000000010000000,
31'b0010100000001000000000001100000,
31'b0001010000000001010100000000000,
31'b1000000100010000000000100001000,
31'b0000010000000000000000000011100,
31'b0010100000000000000000001100000,
31'b0110000001010000000000010000000,
31'b1000000000000000000000001000101,
31'b1000001110000000000000000010000,
31'b0100010000000000001000000000001,
31'b0110000000101000000000010000000,
31'b0111000000000000010000000000100,
31'b0001000000001000001010000000000,
31'b0110000000100010000000010000000,
31'b0110000000100000000000010000000,
31'b0001000000000010001010000000000,
31'b0001000000000000001010000000000,
31'b0010001000000000000010000000000,
31'b0010001000000010000010000000000,
31'b0010001000000100000010000000000,
31'b0000010000000000010000010000000,
31'b0010001000001000000010000000000,
31'b0110000000110000000000010000000,
31'b0010001000001100000010000000000,
31'b0001000000010000001010000000000,
31'b0110000000001010000000010000000,
31'b0110000000001000000000010000000,
31'b1000000101000000000000100001000,
31'b0110000000001100000000010000000,
31'b0110000000000010000000010000000,
31'b0110000000000000000000010000000,
31'b0110000000000110000000010000000,
31'b0110000000000100000000010000000,
31'b0010001000100000000010000000000,
31'b0110000000011000000000010000000,
31'b0101001000000000001000010000000,
31'b0100000000000000000010000000101,
31'b0001010000000000000000000000100,
31'b0110000000010000000000010000000,
31'b0010000000000000011000000000001,
31'b0110000000010100000000010000000,
31'b0110100110000000000000000000000,
31'b1000001000010001010000000000000,
31'b0011000000000000000010100000000,
31'b0001000000000000010100001000000,
31'b1000010000000001000000000000101,
31'b1000011000000000000001000100000,
31'b0011000000001000000010100000000,
31'b0001000011000000001010000000000,
31'b1000010001000000100001000000000,
31'b1000001000000001010000000000000,
31'b0010100000000000010001000000000,
31'b0000000000000000100010000010000,
31'b1000001001000000000100000000100,
31'b1000000000000000100000000000011,
31'b0100100100000000000000000110000,
31'b0000000100000000011000000000010,
31'b0100000000000000001000110000000,
31'b0100100001000000000000000000011,
31'b0000100000000000000000001010000,
31'b0000100000000010000000001010000,
31'b0100110000000000000001000000000,
31'b0110000011000000000000010000000,
31'b0000100000001000000000001010000,
31'b1000110000000000000000000001001,
31'b0100100000000001010000000100000,
31'b0000000000000100010000100000001,
31'b0000100000010000000000001010000,
31'b0000000000000000010000100000001,
31'b0101000000000000000000010101000,
31'b1000001100000100000000000010000,
31'b1000001100000010000000000010000,
31'b1000001100000000000000000010000,
31'b1000010000010000100001000000000,
31'b1000010000000000010100000000001,
31'b0011000001000000000010100000000,
31'b0001000010001000001010000000000,
31'b1000001000010000000100000000100,
31'b0110000010100000000000010000000,
31'b0001000000000001000000001000100,
31'b0001000010000000001010000000000,
31'b1000010000000000100001000000000,
31'b1000010000000010100001000000000,
31'b1000101000000000000000010010000,
31'b0000010010000000010000010000000,
31'b1000001000000000000100000000100,
31'b1000001000000010000100000000100,
31'b1100000000000000100000001010000,
31'b0001010000000000100000001000010,
31'b0100100000000010000000000000011,
31'b0100100000000000000000000000011,
31'b0000100001000000000000001010000,
31'b0100100000000100000000000000011,
31'b0110000010000010000000010000000,
31'b0110000010000000000000010000000,
31'b0001110000000000000010000000010,
31'b1100100000000000000010000010000,
31'b1001001100000000000000000001000,
31'b0100100000010000000000000000011,
31'b0100000000000010000000010110000,
31'b0100000000000000000000010110000,
31'b0010000000000000000101000001000,
31'b0110000010010000000000010000000,
31'b0010000010000000011000000000001,
31'b1110000000000000000100000000001,
31'b0000000000000001000000000001001,
31'b1010000000100000000000000100000,
31'b0010000000000000000001100000100,
31'b1100000000000001000001000000000,
31'b0010000000000000100000011000000,
31'b1010000000101000000000000100000,
31'b0010000000001000000001100000100,
31'b1100000000001001000001000000000,
31'b0010000101000000000010000000000,
31'b1010000000110000000000000100000,
31'b0010000101000100000010000000000,
31'b1100000000010001000001000000000,
31'b0010000101001000000010000000000,
31'b1110000100000000000000001000000,
31'b1100001000000000000100000000010,
31'b1000000010100000000000000010000,
31'b1010000000000010000000000100000,
31'b1010000000000000000000000100000,
31'b1000001000000000000000100001000,
31'b0000100000000000000000000000101,
31'b1010000000001010000000000100000,
31'b1010000000001000000000000100000,
31'b1000001000001000000000100001000,
31'b1000000010010000000000000010000,
31'b1010000000010010000000000100000,
31'b1010000000010000000000000100000,
31'b1000001000010000000000100001000,
31'b1000000010001000000000000010000,
31'b1010001001000000100000000000000,
31'b1000000010000100000000000010000,
31'b1000000010000010000000000010000,
31'b1000000010000000000000000010000,
31'b0010000100010000000010000000000,
31'b1010000001100000000000000100000,
31'b0010000100010100000010000000000,
31'b1100000001000001000001000000000,
31'b0010000100011000000010000000000,
31'b0001000000000101000000000010001,
31'b0000000100000000000000010000101,
31'b0001000000000001000000000010001,
31'b0010000100000000000010000000000,
31'b0010000100000010000010000000000,
31'b0010000100000100000010000000000,
31'b0010010000000000000100100100000,
31'b0010000100001000000010000000000,
31'b0110100000000000100000000100000,
31'b0010000100001100000010000000000,
31'b1100000000000000100000000000101,
31'b1010000001000010000000000100000,
31'b1010000001000000000000000100000,
31'b1001000000000010101000000000000,
31'b1001000000000000101000000000000,
31'b1010001000010000100000000000000,
31'b1010000001001000000000000100000,
31'b0100010100000000010010000000000,
31'b1001000000001000101000000000000,
31'b1001000010000000000000000001000,
31'b1010000001010000000000000100000,
31'b1010000000000000001000100010000,
31'b1001000000010000101000000000000,
31'b1010001000000000100000000000000,
31'b1010001000000010100000000000000,
31'b1010001000000100100000000000000,
31'b1000000011000000000000000010000,
31'b0011000000000000010000000000010,
31'b1010000010100000000000000100000,
31'b0011000000000100010000000000010,
31'b1100000010000001000001000000000,
31'b0101100000000000100000000001000,
31'b1000010100000000000001000100000,
31'b1000000000110010000000000010000,
31'b1000000000110000000000000010000,
31'b1001000001100000000000000001000,
31'b1000000100000001010000000000000,
31'b1000000000101010000000000010000,
31'b1000000000101000000000000010000,
31'b1000000101000000000100000000100,
31'b1000000000100100000000000010000,
31'b1000000000100010000000000010000,
31'b1000000000100000000000000010000,
31'b1010000010000010000000000100000,
31'b1010000010000000000000000100000,
31'b1000001010000000000000100001000,
31'b1000000000011000000000000010000,
31'b1000000001000000001000100100000,
31'b1000000000010100000000000010000,
31'b1000000000010010000000000010000,
31'b1000000000010000000000000010000,
31'b1001000001000000000000000001000,
31'b0000000000000000000010000000011,
31'b1000000000001010000000000010000,
31'b1000000000001000000000000010000,
31'b1000000000000110000000000010000,
31'b1000000000000100000000000010000,
31'b1000000000000010000000000010000,
31'b1000000000000000000000000010000,
31'b1001000000110000000000000001000,
31'b0100100000000100100000000010000,
31'b0110000000000000010011000000000,
31'b0100100000000000100000000010000,
31'b1000000100010000000100000000100,
31'b0000010000000000000100100010000,
31'b0000000100000000000010000110000,
31'b0000000000000000001001000000100,
31'b1001000000100000000000000001000,
31'b1001000000100010000000000001000,
31'b1001000000100100000000000001000,
31'b1001100000000001000000000000100,
31'b1000000100000000000100000000100,
31'b1000000100000010000100000000100,
31'b1000000100000100000100000000100,
31'b1000000001100000000000000010000,
31'b1001000000010000000000000001000,
31'b1010000011000000000000000100000,
31'b1001000000010100000000000001000,
31'b1001000010000000101000000000000,
31'b1000000000000000001000100100000,
31'b1000000001010100000000000010000,
31'b1000000001010010000000000010000,
31'b1000000001010000000000000010000,
31'b1001000000000000000000000001000,
31'b1001000000000010000000000001000,
31'b1001000000000100000000000001000,
31'b1000000001001000000000000010000,
31'b0000010000000000000011000000000,
31'b1000000001000100000000000010000,
31'b1000000001000010000000000010000,
31'b1000000001000000000000000010000,
31'b0010000001010000000010000000000,
31'b1010000100100000000000000100000,
31'b0010000100000000000001100000100,
31'b1100000100000001000001000000000,
31'b0010000100000000100000011000000,
31'b1110000000010000000000001000000,
31'b0000000001000000000000010000101,
31'b0001100000000000000100000001001,
31'b0010000001000000000010000000000,
31'b1000000010000001010000000000000,
31'b0010000001000100000010000000000,
31'b1010010000000000000001000010000,
31'b0010000001001000000010000000000,
31'b1110000000000000000000001000000,
31'b0010000001001100000010000000000,
31'b1110000000000100000000001000000,
31'b1010000100000010000000000100000,
31'b1010000100000000000000000100000,
31'b1000010000000010010000001000000,
31'b1000010000000000010000001000000,
31'b0001010000000000010001000000010,
31'b1100000000000000010001000010000,
31'b0000010010000000000000100000100,
31'b1000010000001000010000001000000,
31'b0010000001100000000010000000000,
31'b1010000100010000000000000100000,
31'b0101000001000000001000010000000,
31'b1000010000010000010000001000000,
31'b0010101000000000000000001100000,
31'b1110000000100000000000001000000,
31'b1000001000000000000000001000101,
31'b1000000110000000000000000010000,
31'b0010000000010000000010000000000,
31'b0010000000010010000010000000000,
31'b0010000000010100000010000000000,
31'b0010010000100000001000000000100,
31'b0010000000011000000010000000000,
31'b0110001000100000000000010000000,
31'b0000000000000000000000010000101,
31'b0001001000000000001010000000000,
31'b0010000000000000000010000000000,
31'b0010000000000010000010000000000,
31'b0010000000000100000010000000000,
31'b0010000000000110000010000000000,
31'b0010000000001000000010000000000,
31'b0100000000000000011000000000100,
31'b0010000000001100000010000000000,
31'b0111010000000000000000000000001,
31'b0010000000110000000010000000000,
31'b0001000000000000010000000000001,
31'b0101000000010000001000010000000,
31'b0010010000000000001000000000100,
31'b0110001000000010000000010000000,
31'b0110001000000000000000010000000,
31'b0100010000000000010010000000000,
31'b0110001000000100000000010000000,
31'b0010000000100000000010000000000,
31'b0010000000100010000010000000000,
31'b0101000000000000001000010000000,
31'b0101000000000010001000010000000,
31'b0010000000101000000010000000000,
31'b0110001000010000000000010000000,
31'b0101000000001000001000010000000,
31'b1000000111000000000000000010000,
31'b1000000001000000000000000100011,
31'b1000000000010001010000000000000,
31'b0011001000000000000010100000000,
31'b1100000000000000000000001110000,
31'b1000010000000010000001000100000,
31'b1000010000000000000001000100000,
31'b0000010000100000000000100000100,
31'b1000010000000100000001000100000,
31'b1000000000000011010000000000000,
31'b1000000000000001010000000000000,
31'b1000100001000000000000010010000,
31'b1000000000000101010000000000000,
31'b1000000001000000000100000000100,
31'b0000000000000000001010100000000,
31'b1000000100100010000000000010000,
31'b1000000100100000000000000010000,
31'b0100100000000000100100000000100,
31'b1010000110000000000000000100000,
31'b0000101000000000000000001010000,
31'b1000010010000000010000001000000,
31'b0000010000000100000000100000100,
31'b1000010000100000000001000100000,
31'b0000010000000000000000100000100,
31'b1000000100010000000000000010000,
31'b1001000101000000000000000001000,
31'b1000000000100001010000000000000,
31'b1000100000000000010000000001100,
31'b1000000100001000000000000010000,
31'b1000000100000110000000000010000,
31'b1000000100000100000000000010000,
31'b1000000100000010000000000010000,
31'b1000000100000000000000000010000,
31'b1000000000000000000000000100011,
31'b1000000001010001010000000000000,
31'b0010100000000000000000000000110,
31'b0100100100000000100000000010000,
31'b1000000000010000000100000000100,
31'b1000010001000000000001000100000,
31'b0000000000000000000010000110000,
31'b0000000100000000001001000000100,
31'b0010000010000000000010000000000,
31'b1000000001000001010000000000000,
31'b1000100000000000000000010010000,
31'b1000100000000010000000010010000,
31'b1000000000000000000100000000100,
31'b1000000000000010000100000000100,
31'b1000000000000100000100000000100,
31'b1000000101100000000000000010000,
31'b1001000100010000000000000001000,
31'b0010000000000001000000000001010,
31'b0010100000100000000000000000110,
31'b0010010010000000001000000000100,
31'b1000000100000000001000100100000,
31'b0110001010000000000000010000000,
31'b0000010001000000000000100000100,
31'b1000010000000000001110000000000,
31'b1001000100000000000000000001000,
31'b1001000100000010000000000001000,
31'b1001000100000100000000000001000,
31'b1001000000000000010100010000000,
31'b1000000000100000000100000000100,
31'b1000000101000100000000000010000,
31'b1000000101000010000000000010000,
31'b1000000101000000000000000010000,
31'b0110110000000000000000000000000,
31'b0110110000000010000000000000000,
31'b1100000001000000110000000000000,
31'b0001000010000000000010010000010,
31'b0110110000001000000000000000000,
31'b1001000000000000000010000100100,
31'b0010000000000000100100100000000,
31'b0001000000010000000100000010000,
31'b0000000001000000000100000001000,
31'b0001100000000000000000010000100,
31'b0000100000101000010000000000000,
31'b0001000000001000000100000010000,
31'b0000100000100100010000000000000,
31'b0001000000000100000100000010000,
31'b0000100000100000010000000000000,
31'b0001000000000000000100000010000,
31'b1010000000000000010100000000010,
31'b1010011000000000000000000100000,
31'b1000010000000000000000100001000,
31'b1000010000000010000000100001000,
31'b0100000001000000000000100000010,
31'b0100100000000000001000010000001,
31'b0000100000010000010000000000000,
31'b0000100000010010010000000000000,
31'b0000100000001100010000000000000,
31'b0001100000100000000000010000100,
31'b0000100000001000010000000000000,
31'b0000100000001010010000000000000,
31'b0000100000000100010000000000000,
31'b0000100000000110010000000000000,
31'b0000100000000000010000000000000,
31'b0000100000000010010000000000000,
31'b0000000000010000000100000001000,
31'b0100000010000000000001010000000,
31'b1100000000000000110000000000000,
31'b0000000100010000010000010000000,
31'b0100000000100000000000100000010,
31'b0100000010001000000001010000000,
31'b1100000000001000110000000000000,
31'b0001010100000000001010000000000,
31'b0000000000000000000100000001000,
31'b0000000000000010000100000001000,
31'b0000000000000100000100000001000,
31'b0000000100000000010000010000000,
31'b0000000000001000000100000001000,
31'b0000000000100001000000010010000,
31'b0000100001100000010000000000000,
31'b0001000001000000000100000010000,
31'b0100000000001000000000100000010,
31'b0100000010100000000001010000000,
31'b1100000000100000110000000000000,
31'b0010001100000000001000000000100,
31'b0100000000000000000000100000010,
31'b0100000000000010000000100000010,
31'b0100000000000100000000100000010,
31'b0100000000000110000000100000010,
31'b0000000000100000000100000001000,
31'b0000000000100010000100000001000,
31'b0000100001001000010000000000000,
31'b0000100000000001000100000000100,
31'b0001000100000000000000000000100,
31'b0000000000000001000000010010000,
31'b0000100001000000010000000000000,
31'b0000100001000010010000000000000,
31'b0110110010000000000000000000000,
31'b0100000001000000000001010000000,
31'b1000000001000000000000010001001,
31'b0001000000000000000010010000010,
31'b1000000100000001000000000000101,
31'b1001000000000000000000010010001,
31'b0010100100000001000000000100000,
31'b0001000010010000000100000010000,
31'b0000100000000000000001001100000,
31'b0110000000000000000000001001100,
31'b0000100010101000010000000000000,
31'b0001000010001000000100000010000,
31'b0000100010100100010000000000000,
31'b0011000000000000000000000000111,
31'b0000100010100000010000000000000,
31'b0001000010000000000100000010000,
31'b0110000000000010001000000000010,
31'b0110000000000000001000000000010,
31'b1000010010000000000000100001000,
31'b0110000000000100001000000000010,
31'b0100100100000000000001000000000,
31'b0110000000001000001000000000010,
31'b0000100010010000010000000000000,
31'b1000100100000000000000000001001,
31'b0000100010001100010000000000000,
31'b1100001000000000000001001000000,
31'b0000100010001000010000000000000,
31'b1000100000000000000000101000100,
31'b0000100010000100010000000000000,
31'b1000100000000000100001010000000,
31'b0000100010000000010000000000000,
31'b1000011000000000000000000010000,
31'b0100000000000010000001010000000,
31'b0100000000000000000001010000000,
31'b1000000000000000000000010001001,
31'b0000000000000000101100000000000,
31'b0100000010100000000000100000010,
31'b0100000000001000000001010000000,
31'b1010000000000001100000001000000,
31'b0000010000000000000000011010000,
31'b0000000010000000000100000001000,
31'b0100000000010000000001010000000,
31'b0000000010000100000100000001000,
31'b0000000110000000010000010000000,
31'b0000001000100000000011000000000,
31'b0100000000011000000001010000000,
31'b0000100011100000010000000000000,
31'b0001000100000000100000001000010,
31'b0100000010001000000000100000010,
31'b0100000000100000000001010000000,
31'b1000010000000000100000000110000,
31'b0010000000000001000000010100000,
31'b0100000010000000000000100000010,
31'b0100000010000010000000100000010,
31'b0101000000000000010001000000100,
31'b1010010000000000001000000001000,
31'b0000001000001000000011000000000,
31'b0100001000000000000000000011010,
31'b0000100011001000010000000000000,
31'b0010100000000000011000100000000,
31'b0000001000000000000011000000000,
31'b0000001000000010000011000000000,
31'b0000100011000000010000000000000,
31'b1010100000000001000010000000000,
31'b0100000001000000001000000000001,
31'b0100100000000000000000110000010,
31'b0100100000000000010000001100000,
31'b0000000001010000010000010000000,
31'b1001000000000000001001000010000,
31'b1000001010000000000001000100000,
31'b0010100010000001000000000100000,
31'b0001010001000000001010000000000,
31'b0000100000000001000000000010000,
31'b0000100000000011000000000010000,
31'b0000100000000101000000000010000,
31'b0000000001000000010000010000000,
31'b0001000001100000000000000000100,
31'b0001000100000100000100000010000,
31'b0000100100100000010000000000000,
31'b0001000100000000000100000010000,
31'b0100100010001000000001000000000,
31'b1000001000000100010000001000000,
31'b1000010100000000000000100001000,
31'b1000001000000000010000001000000,
31'b0100100010000000000001000000000,
31'b0110010001000000000000010000000,
31'b0000100100010000010000000000000,
31'b1000100010000000000000000001001,
31'b0001000001001000000000000000100,
31'b0001000000000001010100000000000,
31'b0000100100001000010000000000000,
31'b0000000000000000000000000011100,
31'b0001000001000000000000000000100,
31'b0001000001000010000000000000100,
31'b0000100100000000010000000000000,
31'b0000100100000010010000000000000,
31'b0100000000000000001000000000001,
31'b0100000000000010001000000000001,
31'b0100000000000100001000000000001,
31'b0000000000010000010000010000000,
31'b0100000000001000001000000000001,
31'b0110010000100000000000010000000,
31'b0100001000100000010010000000000,
31'b0001010000000000001010000000000,
31'b0000000100000000000100000001000,
31'b0000000000000100010000010000000,
31'b0000000000000010010000010000000,
31'b0000000000000000010000010000000,
31'b0001000000100000000000000000100,
31'b0001000000100010000000000000100,
31'b0001000000100100000000000000100,
31'b0000000000001000010000010000000,
31'b0100000000100000001000000000001,
31'b0110010000001000000000010000000,
31'b0100001000001000010010000000000,
31'b0010001000000000001000000000100,
31'b0001000000010000000000000000100,
31'b0110010000000000000000010000000,
31'b0100001000000000010010000000000,
31'b0110010000000100000000010000000,
31'b0001000000001000000000000000100,
31'b0001000000001010000000000000100,
31'b0001000000001100000000000000100,
31'b0000000000100000010000010000000,
31'b0001000000000000000000000000100,
31'b0001000000000010000000000000100,
31'b0001000000000100000000000000100,
31'b0001000000000110000000000000100,
31'b1000000001010000100001000000000,
31'b1000001000001000000001000100000,
31'b0011010000000000000010100000000,
31'b0001010000000000010100001000000,
31'b1000000000000001000000000000101,
31'b1000001000000000000001000100000,
31'b0010100000000001000000000100000,
31'b1000100000100000000000000001001,
31'b1000000001000000100001000000000,
31'b1000011000000001010000000000000,
31'b1010000000000001000010010000000,
31'b0000010000000000100010000010000,
31'b1000000001001000100001000000000,
31'b1000010000000000100000000000011,
31'b0010100000010001000000000100000,
31'b0001000110000000000100000010000,
31'b0100100000001000000001000000000,
31'b0110000100000000001000000000010,
31'b0000110000000000000000001010000,
31'b1000100000001000000000000001001,
31'b0100100000000000000001000000000,
31'b0100100000000010000001000000000,
31'b0000001000000000000000100000100,
31'b1000100000000000000000000001001,
31'b1101000000000001001000000000000,
31'b0011000000000000001000100000100,
31'b0000110000010000000000001010000,
31'b0000010000000000010000100000001,
31'b0100100000010000000001000000000,
31'b0111000000000000000100001000000,
31'b0000100110000000010000000000000,
31'b1000100000010000000000000001001,
31'b1000000000010000100001000000000,
31'b1000000000000000010100000000001,
31'b1000000100000000000000010001001,
31'b0000000100000000101100000000000,
31'b1000000001000001000000000000101,
31'b1000001001000000000001000100000,
31'b0010100001000001000000000100000,
31'b0001010010000000001010000000000,
31'b1000000000000000100001000000000,
31'b1000000000000010100001000000000,
31'b1000000000000100100001000000000,
31'b0000000010000000010000010000000,
31'b1000000000001000100001000000000,
31'b1000000000001010100001000000000,
31'b1000000000001100100001000000000,
31'b0001000000000000100000001000010,
31'b1001100000000000000000000010001,
31'b1000100000000000000011001000000,
31'b0011000000000000000000000110100,
31'b0010001010000000001000000000100,
31'b0100100001000000000001000000000,
31'b0110010010000000000000010000000,
31'b0001100000000000000010000000010,
31'b1000100001000000000000000001001,
31'b1000000000100000100001000000000,
31'b1001000000000000010000101000000,
31'b1001000000000000000000010100010,
31'b0000000010100000010000010000000,
31'b0001000010000000000000000000100,
31'b0001000010000010000000000000100,
31'b0001000010000100000000000000100,
31'b0001000010000110000000000000100,
31'b0010000000000000001100000010000,
31'b1010010000100000000000000100000,
31'b0010010000000000000001100000100,
31'b1100010000000001000001000000000,
31'b1000000000000011000000001010000,
31'b1000000000000001000000001010000,
31'b0010100000000000001000010000100,
31'b1100000000010000010000000100000,
31'b0000100000000000001010000000001,
31'b0001101000000000000000010000100,
31'b0000101000101000010000000000000,
31'b1100000000001000010000000100000,
31'b0000101000100100010000000000000,
31'b1100000000000100010000000100000,
31'b0000101000100000010000000000000,
31'b1100000000000000010000000100000,
31'b1010010000000010000000000100000,
31'b1010010000000000000000000100000,
31'b1000011000000000000000100001000,
31'b1000000100000000010000001000000,
31'b0101100000000000000010000000100,
31'b1010010000001000000000000100000,
31'b0000101000010000010000000000000,
31'b1000010010010000000000000010000,
31'b0000101000001100010000000000000,
31'b1100000010000000000001001000000,
31'b0000101000001000010000000000000,
31'b1000010010001000000000000010000,
31'b0000101000000100010000000000000,
31'b1010000000000001010001000000000,
31'b0000101000000000010000000000000,
31'b1000010010000000000000000010000,
31'b0100000000000001000010000010000,
31'b0100001010000000000001010000000,
31'b1100001000000000110000000000000,
31'b0010000100100000001000000000100,
31'b0100001000100000000000100000010,
31'b0000000010000000000100100010000,
31'b1100000000000001000000000000011,
31'b0011000000000000001100000001000,
31'b0000001000000000000100000001000,
31'b0000001000000010000100000001000,
31'b0000001000000100000100000001000,
31'b0010000000000000000100100100000,
31'b0000001000001000000100000001000,
31'b0000001000100001000000010010000,
31'b0000101001100000010000000000000,
31'b1100000001000000010000000100000,
31'b0100001000001000000000100000010,
31'b1010010001000000000000000100000,
31'b0100000100001000010010000000000,
31'b0010000100000000001000000000100,
31'b0100001000000000000000100000010,
31'b0100001000000010000000100000010,
31'b0100000100000000010010000000000,
31'b0110000000000000000000000101010,
31'b0000001000100000000100000001000,
31'b0100000010000000000000000011010,
31'b0000101001001000010000000000000,
31'b0010000100010000001000000000100,
31'b0000000010000000000011000000000,
31'b0000001000000001000000010010000,
31'b0000101001000000010000000000000,
31'b1000010011000000000000000010000,
31'b0011010000000000010000000000010,
31'b1110000000000000010000000010000,
31'b0001000000000000000100100001000,
31'b0001001000000000000010010000010,
31'b1000000100000010000001000100000,
31'b1000000100000000000001000100000,
31'b0000000100100000000000100000100,
31'b1000010000110000000000000010000,
31'b0000101000000000000001001100000,
31'b1100000000100000000001001000000,
31'b0000000000100000000000001001001,
31'b1010000000000001000000001100000,
31'b0000000001100000000011000000000,
31'b1000010000100100000000000010000,
31'b0000000000000000001100000100000,
31'b1000010000100000000000000010000,
31'b0000000100001100000000100000100,
31'b1100000000010000000001001000000,
31'b0000000100001000000000100000100,
31'b1000010000011000000000000010000,
31'b0000000100000100000000100000100,
31'b1000010000010100000000000010000,
31'b0000000100000000000000100000100,
31'b1000010000010000000000000010000,
31'b0000000001001000000011000000000,
31'b1100000000000000000001001000000,
31'b0000000000000000000000001001001,
31'b1000010000001000000000000010000,
31'b0000000001000000000011000000000,
31'b1000010000000100000000000010000,
31'b0101000000000000000000000000010,
31'b1000010000000000000000000010000,
31'b0100001000000010000001010000000,
31'b0100001000000000000001010000000,
31'b1001100000000000100000000000010,
31'b0000100000000000000000110000100,
31'b0000000000110000000011000000000,
31'b0000000000000000000100100010000,
31'b0000010100000000000010000110000,
31'b0000010000000000001001000000100,
31'b0000001010000000000100000001000,
31'b0100001000010000000001010000000,
31'b0000001010000100000100000001000,
31'b0010100100000001100000000000000,
31'b0000000000100000000011000000000,
31'b0000000000100010000011000000000,
31'b0000000001000000001100000100000,
31'b1000010001100000000000000010000,
31'b0000000000011000000011000000000,
31'b0100001000100000000001010000000,
31'b0010000100000001000010001000000,
31'b0010001000000001000000010100000,
31'b0000000000010000000011000000000,
31'b0000000000100000000100100010000,
31'b0000000101000000000000100000100,
31'b1000010001010000000000000010000,
31'b0000000000001000000011000000000,
31'b0100000000000000000000000011010,
31'b0000000001000000000000001001001,
31'b1001000000000000000010001000010,
31'b0000000000000000000011000000000,
31'b0000000000000010000011000000000,
31'b0000000000000100000011000000000,
31'b1000010001000000000000000010000,
31'b0100100000000000000110000001000,
31'b1000000010001000000001000100000,
31'b1001000000000000100001100000000,
31'b1000000000100000010000001000000,
31'b1001000000000000000000011000100,
31'b1000000010000000000001000100000,
31'b0000000010100000000000100000100,
31'b1000000010000100000001000100000,
31'b0010010001000000000010000000000,
31'b1010000000000100000001000010000,
31'b1010000000000010000001000010000,
31'b1010000000000000000001000010000,
31'b0011000000000000000000001010010,
31'b1110010000000000000000001000000,
31'b0000101100100000010000000000000,
31'b1100000100000000010000000100000,
31'b1000000000000110010000001000000,
31'b1000000000000100010000001000000,
31'b1000000000000010010000001000000,
31'b1000000000000000010000001000000,
31'b0001000000000000010001000000010,
31'b1000000010100000000001000100000,
31'b0000000010000000000000100000100,
31'b1000000000001000010000001000000,
31'b0010010001100000000010000000000,
31'b1100000000000001000000000110000,
31'b1000100000000000000000100010001,
31'b1000000000010000010000001000000,
31'b0001001001000000000000000000100,
31'b0001001001000010000000000000100,
31'b0000101100000000010000000000000,
31'b1000010110000000000000000010000,
31'b0100001000000000001000000000001,
31'b0101000000000000000010010000100,
31'b0100001000000100001000000000001,
31'b0010000000100000001000000000100,
31'b0100001000001000001000000000001,
31'b1000100000000000000100001001000,
31'b0100000000100000010010000000000,
31'b0111000000010000000000000000001,
31'b0010010000000000000010000000000,
31'b0010010000000010000010000000000,
31'b0010010000000100000010000000000,
31'b0000001000000000010000010000000,
31'b0010010000001000000010000000000,
31'b0111000000000100000000000000001,
31'b0111000000000010000000000000001,
31'b0111000000000000000000000000001,
31'b0100001000100000001000000000001,
31'b0010000000000100001000000000100,
31'b0100000000001000010010000000000,
31'b0010000000000000001000000000100,
31'b0100000000000100010010000000000,
31'b0110011000000000000000010000000,
31'b0100000000000000010010000000000,
31'b0100000000000010010010000000000,
31'b0010010000100000000010000000000,
31'b0010010000100010000010000000000,
31'b0101010000000000001000010000000,
31'b0010000000010000001000000000100,
31'b0001001000000000000000000000100,
31'b0001001000000010000000000000100,
31'b0100000000010000010010000000000,
31'b0111000000100000000000000000001,
31'b1000000000001010000001000100000,
31'b1000000000001000000001000100000,
31'b0001000000000000000000001100010,
31'b1000000010100000010000001000000,
31'b1000000000000010000001000100000,
31'b1000000000000000000001000100000,
31'b0000000000100000000000100000100,
31'b1000000000000100000001000100000,
31'b1000010000000011010000000000000,
31'b1000010000000001010000000000000,
31'b0101000000000000001000100000001,
31'b1010000010000000000001000010000,
31'b1000010001000000000100000000100,
31'b1000000000010000000001000100000,
31'b0000000100000000001100000100000,
31'b1000010100100000000000000010000,
31'b0000000000001100000000100000100,
31'b1000000010000100010000001000000,
31'b0000000000001000000000100000100,
31'b1000000010000000010000001000000,
31'b0000000000000100000000100000100,
31'b1000000000100000000001000100000,
31'b0000000000000000000000100000100,
31'b0000000000000010000000100000100,
31'b0010000001000000100000000001100,
31'b1100000100000000000001001000000,
31'b0000000100000000000000001001001,
31'b1000010100001000000000000010000,
31'b0000000101000000000011000000000,
31'b1000010100000100000000000010000,
31'b0000000000010000000000100000100,
31'b1000010100000000000000000010000,
31'b1000010000000000000000000100011,
31'b1000001000000000010100000000001,
31'b0010110000000000000000000000110,
31'b0010100000010001100000000000000,
31'b1000010000010000000100000000100,
31'b1000000001000000000001000100000,
31'b0000010000000000000010000110000,
31'b1000000001000100000001000100000,
31'b1000001000000000100001000000000,
31'b1000010001000001010000000000000,
31'b1000110000000000000000010010000,
31'b0010100000000001100000000000000,
31'b1000010000000000000100000000100,
31'b1000010000000010000100000000100,
31'b1000010000000100000100000000100,
31'b0111000010000000000000000000001,
31'b0010000000010000100000000001100,
31'b0010010000000001000000000001010,
31'b0010000000000001000010001000000,
31'b0010000010000000001000000000100,
31'b0000000100010000000011000000000,
31'b1000000001100000000001000100000,
31'b0000000001000000000000100000100,
31'b1000000000000000001110000000000,
31'b0010000000000000100000000001100,
31'b0100100000000000100001000100000,
31'b0010000000010001000010001000000,
31'b0010100000100001100000000000000,
31'b0000000100000000000011000000000,
31'b0000000100000010000011000000000,
31'b0000000100000100000011000000000,
31'b1000010101000000000000000010000,
31'b0111000000000000000000000000000,
31'b0111000000000010000000000000000,
31'b0111000000000100000000000000000,
31'b0111000000000110000000000000000,
31'b0111000000001000000000000000000,
31'b0111000000001010000000000000000,
31'b0111000000001100000000000000000,
31'b0100001000010000001000000000000,
31'b0111000000010000000000000000000,
31'b0000010000000000000000010000100,
31'b0111000000010100000000000000000,
31'b0100001000001000001000000000000,
31'b0111000000011000000000000000000,
31'b0100001000000100001000000000000,
31'b0100001000000010001000000000000,
31'b0100001000000000001000000000000,
31'b0111000000100000000000000000000,
31'b0111000000100010000000000000000,
31'b0000000000000000001010010000000,
31'b0001001000000000000000000000101,
31'b0111000000101000000000000000000,
31'b1000100001000000000000100010000,
31'b0001010000010000010000000000000,
31'b0110000000000000010000010000100,
31'b0111000000110000000000000000000,
31'b0100000000000000010010000000001,
31'b0001010000001000010000000000000,
31'b0100001000101000001000000000000,
31'b0010000000000000001000000000101,
31'b0100001000100100001000000000000,
31'b0001010000000000010000000000000,
31'b0100001000100000001000000000000,
31'b0111000001000000000000000000000,
31'b0111000001000010000000000000000,
31'b0100000000000000101000000100000,
31'b0110000000001000000000000011000,
31'b1010000000000000000001000010001,
31'b1011000000000000000010001000000,
31'b0110000000000010000000000011000,
31'b0110000000000000000000000011000,
31'b0111000001010000000000000000000,
31'b0100000010000000000000000101000,
31'b1000001000000000001010001000000,
31'b1000001010000001000000000000100,
31'b1000100000000000000111000000000,
31'b0100001001000100001000000000000,
31'b0101000000000000100000100001000,
31'b0100001001000000001000000000000,
31'b0111000001100000000000000000000,
31'b1000100000001000000000100010000,
31'b0001000000000000100100000000010,
31'b1000101000000000101000000000000,
31'b1000100000000010000000100010000,
31'b1000100000000000000000100010000,
31'b0001010001010000010000000000000,
31'b1100000000000000001000011000000,
31'b1000101010000000000000000001000,
31'b0000010000000000010000000011000,
31'b0001010001001000010000000000000,
31'b0010000010000001000001000001000,
31'b1000000000000000010000001000001,
31'b1000100000010000000000100010000,
31'b0001010001000000010000000000000,
31'b0100001001100000001000000000000,
31'b0111000010000000000000000000000,
31'b0111000010000010000000000000000,
31'b0111000010000100000000000000000,
31'b1000010000000000000100000000101,
31'b0100001000000000100000000001000,
31'b0101000001000000001000100000000,
31'b1000001000010000010100000000000,
31'b1000010000010000000000000100010,
31'b0111000010010000000000000000000,
31'b0100000001000000000000000101000,
31'b1000001000001000010100000000000,
31'b1000010000001000000000000100010,
31'b1000001000000100010100000000000,
31'b1000010000000100000000000100010,
31'b1000001000000000010100000000000,
31'b1000010000000000000000000100010,
31'b1100000100000000000010000001000,
31'b0000000101001000000000001001000,
31'b0001000100000000000000001010000,
31'b0000000100000000000011000000001,
31'b0101010100000000000001000000000,
31'b0000000101000000000000001001000,
31'b0001010010010000010000000000000,
31'b0010000001000000000010110000000,
31'b1000101001000000000000000001000,
31'b0000000001000000000000100000101,
31'b0001010010001000010000000000000,
31'b0010000100000000100000101000000,
31'b0011000000000001000001000010000,
31'b0010000100000000000001010000100,
31'b0001010010000000010000000000000,
31'b1001101000000000000000000010000,
31'b0111000011000000000000000000000,
31'b0100000000010000000000000101000,
31'b1000011000000000100000000000010,
31'b1000001000010001000000000000100,
31'b0101000000000010001000100000000,
31'b0101000000000000001000100000000,
31'b1000010000000001010000000000001,
31'b0110000010000000000000000011000,
31'b0100000000000010000000000101000,
31'b0100000000000000000000000101000,
31'b1000000000000000000001000100001,
31'b1000001000000001000000000000100,
31'b0110000000000000101000000010000,
31'b0100000000001000000000000101000,
31'b1000001001000000010100000000000,
31'b1000010001000000000000000100010,
31'b1000101000010000000000000001000,
31'b0000000100001000000000001001000,
31'b0001000101000000000000001010000,
31'b0010000000010001000001000001000,
31'b0000011000000000010000100000000,
31'b0000000100000000000000001001000,
31'b0000010100000000000010000000010,
31'b0010000000000000000010110000000,
31'b1000101000000000000000000001000,
31'b0000000000000000000000100000101,
31'b1000101000000100000000000001000,
31'b0010000000000001000001000001000,
31'b1000101000001000000000000001000,
31'b0000000100010000000000001001000,
31'b0001010011000000010000000000000,
31'b0010000000010000000010110000000,
31'b1000000000000000000000110010000,
31'b1100000000010001000000000000010,
31'b1100100000000000001000001000000,
31'b0000100010000000010100001000000,
31'b1100001000000000000101000000000,
31'b0000100001000100001010000000000,
31'b1000100000000000000100100000100,
31'b0000100001000000001010000000000,
31'b0010000000000000000000100000110,
31'b1100000000000001000000000000010,
31'b0011000010000000010001000000000,
31'b1100000000000101000000000000010,
31'b0011000000100000000000001100000,
31'b1100000000001001000000000000010,
31'b0101000000000001000001001000000,
31'b0100001100000000001000000000000,
31'b1100000010000000000010000001000,
31'b0000101001000000010000000000001,
31'b0001000010000000000000001010000,
31'b0000001000000000001000001100000,
31'b0110000000000000000100000001100,
31'b0000100000000000000101000100000,
31'b0001010100010000010000000000000,
31'b0000100001100000001010000000000,
31'b0011000000001000000000001100000,
31'b1100000000100001000000000000010,
31'b0001010100001000010000000000000,
31'b1100000000000000101010000000000,
31'b0011000000000000000000001100000,
31'b0011000000000010000000001100000,
31'b0001010100000000010000000000000,
31'b0100001100100000001000000000000,
31'b1100000000000000010000000100001,
31'b0000101000100000010000000000001,
31'b0110100000000000010000000000100,
31'b0000100000001000001010000000000,
31'b0000110000110000000000000000100,
31'b0000100000000100001010000000000,
31'b0000100000000010001010000000000,
31'b0000100000000000001010000000000,
31'b0011101000000000000010000000000,
31'b1100000001000001000000000000010,
31'b1000000000000010001000010100000,
31'b1000000000000000001000010100000,
31'b0000110000100000000000000000100,
31'b0000010000000101000000000001000,
31'b0000010000000011000000000001000,
31'b0000010000000001000000000001000,
31'b1000010010000000000000000010001,
31'b0000101000000000010000000000001,
31'b0001000100000000100100000000010,
31'b0000101000000100010000000000001,
31'b0000110000010000000000000000100,
31'b0000000010000000000000001001000,
31'b0000010010000000000010000000010,
31'b0000100000100000001010000000000,
31'b0000110000001000000000000000100,
31'b0000110000001010000000000000100,
31'b0000010000000000000100010010000,
31'b1010000000000001100100000000000,
31'b0000110000000000000000000000100,
31'b0000110000000010000000000000100,
31'b0000000000000000101000001000000,
31'b0000010000100001000000000001000,
31'b1100000000100000000010000001000,
31'b0000101000000000000010000101000,
31'b0010100000000000000010100000000,
31'b0000100000000000010100001000000,
31'b0101010000100000000001000000000,
31'b0000001000000000011001000000000,
31'b0011010000000001000000000100000,
31'b0000100011000000001010000000000,
31'b0011000000000100010001000000000,
31'b1100000010000001000000000000010,
31'b0011000000000000010001000000000,
31'b0011000000000010010001000000000,
31'b1000001000000010000000010001000,
31'b1000001000000000000000010001000,
31'b1010000000000000000000110100000,
31'b1000010100000000000000000100010,
31'b1100000000000000000010000001000,
31'b0000000001001000000000001001000,
31'b0001000000000000000000001010000,
31'b0000000000000000000011000000001,
31'b0101010000000000000001000000000,
31'b0000000001000000000000001001000,
31'b0001000000001000000000001010000,
31'b0000000001000100000000001001000,
31'b1100000000010000000010000001000,
31'b0010000000001000000001010000100,
31'b0001000000010000000000001010000,
31'b0010000000000000100000101000000,
31'b0101010000010000000001000000000,
31'b0010000000000000000001010000100,
31'b0001010110000000010000000000000,
31'b0010000000001000100000101000000,
31'b1000010000100000000000000010001,
31'b0000000000101000000000001001000,
31'b0011001000000000000000000000110,
31'b0000100010001000001010000000000,
31'b0000010000000001101000000000000,
31'b0000000000100000000000001001000,
31'b0000100000000001000000001000100,
31'b0000100010000000001010000000000,
31'b0110000000000000010010000000010,
31'b0100000100000000000000000101000,
31'b1001001000000000000000010010000,
31'b1000001100000001000000000000100,
31'b0000100000000000100010000001000,
31'b0000000000000000001000000000110,
31'b0000100000010001000000001000100,
31'b0000010010000001000000000001000,
31'b1000010000000000000000000010001,
31'b0000000000001000000000001001000,
31'b0001000001000000000000001010000,
31'b0000000001000000000011000000001,
31'b0000000000000010000000001001000,
31'b0000000000000000000000001001000,
31'b0000010000000000000010000000010,
31'b0000000000000100000000001001000,
31'b1000101100000000000000000001000,
31'b0000000100000000000000100000101,
31'b0001000001010000000000001010000,
31'b0010000100000001000001000001000,
31'b0000110010000000000000000000100,
31'b0000000000010000000000001001000,
31'b0000010000010000000010000000010,
31'b0000000000010100000000001001000,
31'b0111001000000000000000000000000,
31'b0111001000000010000000000000000,
31'b0111001000000100000000000000000,
31'b0100000000011000001000000000000,
31'b0000000000000000010000010000001,
31'b0100000000010100001000000000000,
31'b0100000000010010001000000000000,
31'b0100000000010000001000000000000,
31'b0111001000010000000000000000000,
31'b0100000000001100001000000000000,
31'b0100000000001010001000000000000,
31'b0100000000001000001000000000000,
31'b0100000000000110001000000000000,
31'b0100000000000100001000000000000,
31'b0100000000000010001000000000000,
31'b0100000000000000001000000000000,
31'b0111001000100000000000000000000,
31'b0010010000000000011000000000000,
31'b0001000000000010000000000000101,
31'b0001000000000000000000000000101,
31'b0100010000000000000010000000100,
31'b0100010000000010000010000000100,
31'b0100010000000100000010000000100,
31'b0100000000110000001000000000000,
31'b1000100011000000000000000001000,
31'b0100001000000000010010000000001,
31'b0110010000000000000000010000001,
31'b0100000000101000001000000000000,
31'b0100010000010000000010000000100,
31'b0100000000100100001000000000000,
31'b0100000000100010001000000000000,
31'b0100000000100000001000000000000,
31'b0111001001000000000000000000000,
31'b1000100000000001000010000000010,
31'b1000010010000000100000000000010,
31'b1000100000100000101000000000000,
31'b0100000000000000000000100110000,
31'b0100000001010100001000000000000,
31'b0100000001010010001000000000000,
31'b0100000001010000001000000000000,
31'b1000100010100000000000000001000,
31'b1000010000000000001000000001010,
31'b1000000000000000001010001000000,
31'b1000000010000001000000000000100,
31'b0100000001000110001000000000000,
31'b0100000001000100001000000000000,
31'b0100000001000010001000000000000,
31'b0100000001000000001000000000000,
31'b1000100010010000000000000001000,
31'b1000010000000000000000001000100,
31'b1000100000000010101000000000000,
31'b1000100000000000101000000000000,
31'b0000010010000000010000100000000,
31'b1000101000000000000000100010000,
31'b0010000010000000000100000001010,
31'b1100000000000000000001000010100,
31'b1000100010000000000000000001000,
31'b1000100010000010000000000001000,
31'b1000100010000100000000000001000,
31'b1000100000010000101000000000000,
31'b1000100010001000000000000001000,
31'b0100000001100100001000000000000,
31'b0100010100000000000001100000000,
31'b0100000001100000001000000000000,
31'b0100000000001000100000000001000,
31'b0110000000000000001000000110000,
31'b1000010001000000100000000000010,
31'b1000000001010001000000000000100,
31'b0100000000000000100000000001000,
31'b0100000000000010100000000001000,
31'b1000000000010000010100000000000,
31'b1000000000000000100001000000001,
31'b1000100001100000000000000001000,
31'b1000000100001000000000010001000,
31'b1000000000001000010100000000000,
31'b1000000001000001000000000000100,
31'b1000000000000100010100000000000,
31'b1000000100000000000000010001000,
31'b1000000000000000010100000000000,
31'b0100000010000000001000000000000,
31'b1110010000000000000100000000000,
31'b0011000000000000000100000010010,
31'b0001001100000000000000001010000,
31'b0001000010000000000000000000101,
31'b0100000000100000100000000001000,
31'b0100010000000001001000001000000,
31'b1010100000000000100000100000000,
31'b1001100000010000000000000010000,
31'b1000100001000000000000000001000,
31'b1001000000000000000100010000100,
31'b1000100001000100000000000001000,
31'b1001100000001000000000000010000,
31'b1000100001001000000000000001000,
31'b1001100000000100000000000010000,
31'b1000000000100000010100000000000,
31'b1001100000000000000000000010000,
31'b1000100000110000000000000001000,
31'b1000000000010101000000000000100,
31'b1000010000000000100000000000010,
31'b1000000000010001000000000000100,
31'b0100000001000000100000000001000,
31'b0101001000000000001000100000000,
31'b1000010000001000100000000000010,
31'b1000000001000000100001000000001,
31'b1000100000100000000000000001000,
31'b1000000000000101000000000000100,
31'b0110000000000000000000100000000,
31'b1000000000000001000000000000100,
31'b1000100000101000000000000001000,
31'b1000000101000000000000010001000,
31'b1000000001000000010100000000000,
31'b1000000000001001000000000000100,
31'b1000100000010000000000000001000,
31'b1000100000010010000000000001000,
31'b1000100000010100000000000001000,
31'b1000100010000000101000000000000,
31'b0000010000000000010000100000000,
31'b0000010000000010010000100000000,
31'b0010000000000000000100000001010,
31'b0010001000000000000010110000000,
31'b1000100000000000000000000001000,
31'b1000100000000010000000000001000,
31'b1000100000000100000000000001000,
31'b1000000000100001000000000000100,
31'b1000100000001000000000000001000,
31'b1000100000001010000000000001000,
31'b1000100000001100000000000001000,
31'b1001100001000000000000000010000,
31'b1100000000001000000101000000000,
31'b0000100010000000000010000101000,
31'b1000010000000000000100001010000,
31'b0000000000100000001000001100000,
31'b1100000000000000000101000000000,
31'b0000000010000000011001000000000,
31'b1000000000000000101000010000000,
31'b0000000000000000000100000001001,
31'b0011100001000000000010000000000,
31'b1100001000000001000000000000010,
31'b0110100000000000000001000000010,
31'b0100000100001000001000000000000,
31'b1100000000010000000101000000000,
31'b1000000010000000000000010001000,
31'b0100000100000010001000000000000,
31'b0100000100000000001000000000000,
31'b0000100001000010010000000000001,
31'b0000100001000000010000000000001,
31'b0000000000000010001000001100000,
31'b0000000000000000001000001100000,
31'b1100000000100000000101000000000,
31'b0000101000000000000101000100000,
31'b1010000000000001000100000100000,
31'b0000000000100000000100000001001,
31'b0000100000000001000000000100010,
31'b0100000000000100000000100000011,
31'b0100100001000000001000010000000,
31'b0100000000000000000000100000011,
31'b0011001000000000000000001100000,
31'b1100000000000000000010100010000,
31'b0100010001000000000001100000000,
31'b0100000100100000001000000000000,
31'b0010000000000000010001100000000,
31'b0000100000100000010000000000001,
31'b0011000010000000000000000000110,
31'b0000101000001000001010000000000,
31'b1100000001000000000101000000000,
31'b0000101000000100001010000000000,
31'b1001000000000000000110000000010,
31'b0000101000000000001010000000000,
31'b0011100000000000000010000000000,
31'b0011100000000010000010000000000,
31'b1001000010000000000000010010000,
31'b1000001000000000001000010100000,
31'b0011100000001000000010000000000,
31'b1100010000000000000000000100100,
31'b0100010000100000000001100000000,
31'b0100000101000000001000000000000,
31'b0000100000000010010000000000001,
31'b0000100000000000010000000000001,
31'b0100100000010000001000010000000,
31'b0000100000000100010000000000001,
31'b0000111000010000000000000000100,
31'b0000100000001000010000000000001,
31'b1100000000000000001010000100000,
31'b0000101000100000001010000000000,
31'b0000000000000000000000101010000,
31'b0000100000010000010000000000001,
31'b0100100000000000001000010000000,
31'b0100100000000010001000010000000,
31'b0000111000000000000000000000100,
31'b1000010000000000000000100001001,
31'b0100010000000000000001100000000,
31'b0100010000000010000001100000000,
31'b0110000000000000000011000000100,
31'b0000100000000000000010000101000,
31'b0011000001000000000000000000110,
31'b0000101000000000010100001000000,
31'b0100000100000000100000000001000,
31'b0000000000000000011001000000000,
31'b1000000100010000010100000000000,
31'b0000000010000000000100000001001,
31'b1000000000100001000100000010000,
31'b1000000000001000000000010001000,
31'b1001000001000000000000010010000,
31'b1000000101000001000000000000100,
31'b1000000000000010000000010001000,
31'b1000000000000000000000010001000,
31'b1000000100000000010100000000000,
31'b1000000000000100000000010001000,
31'b1100001000000000000010000001000,
31'b0000100011000000010000000000001,
31'b0001001000000000000000001010000,
31'b0000001000000000000011000000001,
31'b0101011000000000000001000000000,
31'b0000001001000000000000001001000,
31'b0010100000000001000000000010010,
31'b0000001001000100000000001001000,
31'b1000000000000001000100000010000,
31'b1000000000101000000000010001000,
31'b1001000000000000010000000001100,
31'b0110010000000000001001000000000,
31'b1000000000100010000000010001000,
31'b1000000000100000000000010001000,
31'b1000100000000001000000010000100,
31'b1001100100000000000000000010000,
31'b0011000000000100000000000000110,
31'b0000100010100000010000000000001,
31'b0011000000000000000000000000110,
31'b1010000000000000100000110000000,
31'b0100000101000000100000000001000,
31'b0000001000100000000000001001000,
31'b0011000000001000000000000000110,
31'b0000101010000000001010000000000,
31'b1001000000000100000000010010000,
31'b1000000100000101000000000000100,
31'b1001000000000000000000010010000,
31'b1000000100000001000000000000100,
31'b1001100000000000000100000000100,
31'b1000000001000000000000010001000,
31'b1001000000001000000000010010000,
31'b1000000100001001000000000000100,
31'b1000100100010000000000000001000,
31'b0000100010000000010000000000001,
31'b0011000000100000000000000000110,
31'b0000100010000100010000000000001,
31'b0000010100000000010000100000000,
31'b0000001000000000000000001001000,
31'b0010000000000000000000101100000,
31'b0000001000000100000000001001000,
31'b1000100100000000000000000001000,
31'b1000100100000010000000000001000,
31'b1001000000100000000000010010000,
31'b1000100000000000010100010000000,
31'b1000100100001000000000000001000,
31'b1000000000000000010000000010100,
31'b0110000000000000001000000000011,
31'b1001000000000001000100000001000,
31'b0111010000000000000000000000000,
31'b0000000000010000000000010000100,
31'b0111010000000100000000000000000,
31'b0010000000001000000010000000001,
31'b0111010000001000000000000000000,
31'b0010000000000100000010000000001,
31'b0010000000000010000010000000001,
31'b0010000000000000000010000000001,
31'b0000000000000010000000010000100,
31'b0000000000000000000000010000100,
31'b0001000000101000010000000000000,
31'b0000000000000100000000010000100,
31'b0001000000100100010000000000000,
31'b0000000000001000000000010000100,
31'b0001000000100000010000000000000,
31'b0000100000000000000100000010000,
31'b0111010000100000000000000000000,
31'b0010001000000000011000000000000,
31'b0001000000011000010000000000000,
31'b0010001000000100011000000000000,
31'b0100001000000000000010000000100,
31'b0101000000000000001000010000001,
31'b0001000000010000010000000000000,
31'b0010000000100000000010000000001,
31'b0001000000001100010000000000000,
31'b0000000000100000000000010000100,
31'b0001000000001000010000000000000,
31'b0001000000001010010000000000000,
31'b0001000000000100010000000000000,
31'b0001000000000110010000000000000,
31'b0001000000000000010000000000000,
31'b0001000000000010010000000000000,
31'b0111010001000000000000000000000,
31'b0010000000000000000001001001000,
31'b1110000000000000000000001000001,
31'b0010000001001000000010000000001,
31'b0000100100110000000000000000100,
31'b0010000001000100000010000000001,
31'b1011000000000000000000000001010,
31'b0010000001000000000010000000001,
31'b0001100000000000000100000001000,
31'b0000000001000000000000010000100,
31'b0001100000000100000100000001000,
31'b0000000100001001000000000001000,
31'b0000100100100000000000000000100,
31'b0000000100000101000000000001000,
31'b0001000001100000010000000000000,
31'b0000000100000001000000000001000,
31'b1000001000000010000000001000100,
31'b1000001000000000000000001000100,
31'b0001010000000000100100000000010,
31'b1100000000000000100100000010000,
31'b0000100100010000000000000000100,
31'b1000110000000000000000100010000,
31'b0001000001010000010000000000000,
31'b0010000010000000010000000101000,
31'b0000100100001000000000000000100,
31'b0000000000000000010000000011000,
31'b0001000001001000010000000000000,
31'b0001000000000001000100000000100,
31'b0000100100000000000000000000100,
31'b0000100100000010000000000000100,
31'b0001000001000000010000000000000,
31'b0001000001000010010000000000000,
31'b0111010010000000000000000000000,
31'b0010100000000000000100000100000,
31'b1000001001000000100000000000010,
31'b1000000000000000000100000000101,
31'b0101000100100000000001000000000,
31'b1000100000000000000000010010001,
31'b1000000001000001010000000000001,
31'b1000000000010000000000000100010,
31'b0001000000000000000001001100000,
31'b0000000010000000000000010000100,
31'b1000000000001010000000000100010,
31'b1000000000001000000000000100010,
31'b1000000000000110000000000100010,
31'b1000000000000100000000000100010,
31'b1000000000000010000000000100010,
31'b1000000000000000000000000100010,
31'b1110001000000000000100000000000,
31'b0010100000100000000100000100000,
31'b0001010100000000000000001010000,
31'b1100000100000000000000001000010,
31'b0101000100000000000001000000000,
31'b0101000100000010000001000000000,
31'b0001000010010000010000000000000,
31'b1001000100000000000000000001001,
31'b0001000010001100010000000000000,
31'b0000000010100000000000010000100,
31'b0001000010001000010000000000000,
31'b1001000000000000000000101000100,
31'b0001000010000100010000000000000,
31'b1001000000000000100001010000000,
31'b0001000010000000010000000000000,
31'b1000000000100000000000000100010,
31'b1000001000000100100000000000010,
31'b0101100000000000000001010000000,
31'b1000001000000000100000000000010,
31'b1000001000000010100000000000010,
31'b0000001000100000010000100000000,
31'b0101010000000000001000100000000,
31'b1000000000000001010000000000001,
31'b1000000001010000000000000100010,
31'b0110000000000000000100011000000,
31'b0100010000000000000000000101000,
31'b1000010000000000000001000100001,
31'b1000011000000001000000000000100,
31'b0010101000000000100100000000000,
31'b1100000000000001001000010000000,
31'b1000000001000010000000000100010,
31'b1000000001000000000000000100010,
31'b1000000100000000000000000010001,
31'b1000001010000000000000001000100,
31'b0000000100001000000010000000010,
31'b0100100000000000100000000100010,
31'b0000001000000000010000100000000,
31'b0000010100000000000000001001000,
31'b0000000100000000000010000000010,
31'b0010000000000000010000000101000,
31'b1000111000000000000000000001000,
31'b0000010000000000000000100000101,
31'b0001000011001000010000000000000,
31'b0011000000000000011000100000000,
31'b0000100110000000000000000000100,
31'b0000101000000000000000001010001,
31'b0001000011000000010000000000000,
31'b1011000000000001000010000000000,
31'b1100000000000000100000000000100,
31'b0010000000000001100000100000000,
31'b1100000000000100100000000000100,
31'b0010000100001000000010000000001,
31'b1100000000001000100000000000100,
31'b0010000100000100000010000000001,
31'b0011000010000001000000000100000,
31'b0010000100000000000010000000001,
31'b0001000000000001000000000010000,
31'b0000000100000000000000010000100,
31'b0001000000000101000000000010000,
31'b0000000100000100000000010000100,
31'b0001000000001001000000000010000,
31'b0000000100001000000000010000100,
31'b0001000100100000010000000000000,
31'b0000000001000001000000000001000,
31'b1100000000100000100000000000100,
31'b0010001100000000011000000000000,
31'b0001010010000000000000001010000,
31'b1100000010000000000000001000010,
31'b0101000010000000000001000000000,
31'b0101000010000010000001000000000,
31'b0001000100010000010000000000000,
31'b1010000000000001010000000000010,
31'b0001000000100001000000000010000,
31'b0000100000000001010100000000000,
31'b0001000100001000010000000000000,
31'b0001100000000000000000000011100,
31'b0000100001000000000000000000100,
31'b0001000000000000000100010001000,
31'b0001000100000000010000000000000,
31'b0001000100000010010000000000000,
31'b1100000001000000100000000000100,
31'b0010000100000000000001001001000,
31'b0000001010000001000000100010000,
31'b0000000000011001000000000001000,
31'b0000100000110000000000000000100,
31'b0000000000010101000000000001000,
31'b0000000010100000000010000000010,
31'b0000000000010001000000000001000,
31'b0001000001000001000000000010000,
31'b0000000101000000000000010000100,
31'b0000000000100000000100010010000,
31'b0000000000001001000000000001000,
31'b0000100000100000000000000000100,
31'b0000000000000101000000000001000,
31'b0000000000000011000000000001000,
31'b0000000000000001000000000001000,
31'b1000000010000000000000000010001,
31'b1000001100000000000000001000100,
31'b0000000010001000000010000000010,
31'b0100000010000000000001000011000,
31'b0000100000010000000000000000100,
31'b0000100000010010000000000000100,
31'b0000000010000000000010000000010,
31'b0000000010000010000010000000010,
31'b0000100000001000000000000000100,
31'b0000100000001010000000000000100,
31'b0000000000000000000100010010000,
31'b0000000000101001000000000001000,
31'b0000100000000000000000000000100,
31'b0000100000000010000000000000100,
31'b0000100000000100000000000000100,
31'b0000000000100001000000000001000,
31'b1100000010000000100000000000100,
31'b0010100100000000000100000100000,
31'b0011000000001001000000000100000,
31'b1100000000100000000000001000010,
31'b0101000000100000000001000000000,
31'b0101000000100010000001000000000,
31'b0011000000000001000000000100000,
31'b1001000000100000000000000001001,
31'b0001000010000001000000000010000,
31'b0000001000000001001000000100000,
31'b0011010000000000010001000000000,
31'b1100000000000000001000000001100,
31'b0101000000110000000001000000000,
31'b1000011000000000000000010001000,
31'b1010000000000000010010000001000,
31'b1000000100000000000000000100010,
31'b1000000001000000000000000010001,
31'b1100000000000100000000001000010,
31'b0001010000000000000000001010000,
31'b1100000000000000000000001000010,
31'b0101000000000000000001000000000,
31'b0101000000000010000001000000000,
31'b0000000001000000000010000000010,
31'b1001000000000000000000000001001,
31'b1100100000000001001000000000000,
31'b0010100000000000001000100000100,
31'b0001010000010000000000001010000,
31'b1100000000010000000000001000010,
31'b0101000000010000000001000000000,
31'b0110100000000000000100001000000,
31'b0001000110000000010000000000000,
31'b1001000000010000000000000001001,
31'b1000000000100000000000000010001,
31'b1010000000000000100100001000000,
31'b0000001000000001000000100010000,
31'b0100001000010000000000010000010,
31'b0000000000000001101000000000000,
31'b0000010000100000000000001001000,
31'b0000000000100000000010000000010,
31'b0000000010010001000000000001000,
31'b1001100000000000100001000000000,
31'b0100010100000000000000000101000,
31'b0100001000000010000000010000010,
31'b0100001000000000000000010000010,
31'b0000100010100000000000000000100,
31'b0000010000000000001000000000110,
31'b0000000010000011000000000001000,
31'b0000000010000001000000000001000,
31'b1000000000000000000000000010001,
31'b1000000000000010000000000010001,
31'b0000000000001000000010000000010,
31'b0100000000000000000001000011000,
31'b0000000000000100000010000000010,
31'b0000010000000000000000001001000,
31'b0000000000000000000010000000010,
31'b0000000000000010000010000000010,
31'b1000000000010000000000000010001,
31'b1000100000000000010000101000000,
31'b0000000010000000000100010010000,
31'b0100001000100000000000010000010,
31'b0000100010000000000000000000100,
31'b0000100010000010000000000000100,
31'b0000000000010000000010000000010,
31'b0000000010100001000000000001000,
31'b0111011000000000000000000000000,
31'b0010000000100000011000000000000,
31'b1000000100000000000100001010000,
31'b0101000000000000010010010000000,
31'b0100000000100000000010000000100,
31'b0100010000010100001000000000000,
31'b0100010000010010001000000000000,
31'b0100010000010000001000000000000,
31'b0001000000000000001010000000001,
31'b0000001000000000000000010000100,
31'b0110000000100000000000010000001,
31'b0100010000001000001000000000000,
31'b0100010000000110001000000000000,
31'b0100010000000100001000000000000,
31'b0100010000000010001000000000000,
31'b0100010000000000001000000000000,
31'b0100000000001000000010000000100,
31'b0010000000000000011000000000000,
31'b0110000000010000000000010000001,
31'b0010000000000100011000000000000,
31'b0100000000000000000010000000100,
31'b0100000000000010000010000000100,
31'b0100000000000100000010000000100,
31'b0100010000110000001000000000000,
31'b0110000000000100000000010000001,
31'b0010000000010000011000000000000,
31'b0110000000000000000000010000001,
31'b0110000000000010000000010000001,
31'b0100000000010000000010000000100,
31'b0100010000100100001000000000000,
31'b0001001000000000010000000000000,
31'b0100010000100000001000000000000,
31'b1000000010000100100000000000010,
31'b1000000000100000000000001000100,
31'b1000000010000000100000000000010,
31'b1000000010000010100000000000010,
31'b0000000010100000010000100000000,
31'b1001000000000000000000100100010,
31'b1001000000000000010000011000000,
31'b0100010001010000001000000000000,
31'b1000100000000000100010000000100,
31'b1000000000000000001000000001010,
31'b1000010000000000001010001000000,
31'b1000010010000001000000000000100,
31'b0010100010000000100100000000000,
31'b1100000100000000000000000100100,
31'b0100010001000010001000000000000,
31'b0100010001000000001000000000000,
31'b1000000000000010000000001000100,
31'b1000000000000000000000001000100,
31'b1000000010100000100000000000010,
31'b1000000000000100000000001000100,
31'b0000000010000000010000100000000,
31'b1000000000001000000000001000100,
31'b0001000000000000000001000000110,
31'b1000000000001100000000001000100,
31'b1000110010000000000000000001000,
31'b1000000000010000000000001000100,
31'b0110000001000000000000010000001,
31'b1000000000010100000000001000100,
31'b0000101100000000000000000000100,
31'b1000000100000000000000100001001,
31'b0100000100000000000001100000000,
31'b0100010001100000001000000000000,
31'b1110000000100000000100000000000,
31'b0010101000000000000100000100000,
31'b1000000001000000100000000000010,
31'b1000001000000000000100000000101,
31'b0100010000000000100000000001000,
31'b0100010000000010100000000001000,
31'b1000010000010000010100000000000,
31'b1000010000000000100001000000001,
31'b0001001000000000000001001100000,
31'b0000001010000000000000010000100,
31'b1000010000001000010100000000000,
31'b1000010001000001000000000000100,
31'b1010000000000000000000100001010,
31'b1000010100000000000000010001000,
31'b1000010000000000010100000000000,
31'b1000001000000000000000000100010,
31'b1110000000000000000100000000000,
31'b0010000010000000011000000000000,
31'b1110000000000100000100000000000,
31'b0010000010000100011000000000000,
31'b0000000001000000010000100000000,
31'b0100000000000001001000001000000,
31'b0100100000010000000000000000010,
31'b0100100000010010000000000000010,
31'b1110000000010000000100000000000,
31'b0010000100000000100100010000000,
31'b0100100000001000000000000000010,
31'b0110000100000000001001000000000,
31'b0100100000000100000000000000010,
31'b0100100000000110000000000000010,
31'b0100100000000000000000000000010,
31'b0100100000000010000000000000010,
31'b1000000000000100100000000000010,
31'b1000000010100000000000001000100,
31'b1000000000000000100000000000010,
31'b1000000000000010100000000000010,
31'b0000000000100000010000100000000,
31'b0001000000000000100001001000000,
31'b1000000000001000100000000000010,
31'b1000000000001010100000000000010,
31'b1000110000100000000000000001000,
31'b1000010000000101000000000000100,
31'b1000000000010000100000000000010,
31'b1000010000000001000000000000100,
31'b0010100000000000100100000000000,
31'b0011000000000000000010100000001,
31'b1000010001000000010100000000000,
31'b1000010000001001000000000000100,
31'b0000000000001000010000100000000,
31'b1000000010000000000000001000100,
31'b1000000000100000100000000000010,
31'b1000000010000100000000001000100,
31'b0000000000000000010000100000000,
31'b0000000000000010010000100000000,
31'b0000000000000100010000100000000,
31'b0000000000000110010000100000000,
31'b1000110000000000000000000001000,
31'b1000110000000010000000000001000,
31'b1000110000000100000000000001000,
31'b1000100000000000000010001000010,
31'b0000000000010000010000100000000,
31'b0000100000000000000000001010001,
31'b0100100001000000000000000000010,
31'b0100100001000010000000000000010,
31'b1100001000000000100000000000100,
31'b0010001000000001100000100000000,
31'b1000000000000000000100001010000,
31'b1010000000100000100000000000001,
31'b1100010000000000000101000000000,
31'b0010000000000101001000000010000,
31'b1000010000000000101000010000000,
31'b0010000000000001001000000010000,
31'b0001001000000001000000000010000,
31'b0000001100000000000000010000100,
31'b1001000000000000110010000000000,
31'b0100010100001000001000000000000,
31'b0010100000000000000000001010010,
31'b1100000001000000000000000100100,
31'b0100010100000010001000000000000,
31'b0100010100000000001000000000000,
31'b0110000000000000100001000001000,
31'b0010000100000000011000000000000,
31'b1010000000000010100000000000001,
31'b1010000000000000100000000000001,
31'b0100000100000000000010000000100,
31'b0100000100000010000010000000100,
31'b0100000100000100000010000000100,
31'b1010000000001000100000000000001,
31'b0001001000100001000000000010000,
31'b0010000100010000011000000000000,
31'b1010000000000000010101000000000,
31'b1010000000010000100000000000001,
31'b0001000000000000000010100000010,
31'b1000000001000000000000100001001,
31'b0100000001000000000001100000000,
31'b0100010100100000001000000000000,
31'b0011000000000001001000000001000,
31'b1100000000000000000100000000011,
31'b0000000010000001000000100010000,
31'b0100000010010000000000010000010,
31'b0010100000000000011000010000000,
31'b1100000000010000000000000100100,
31'b0100000000110000000001100000000,
31'b0100000000000000000110000010000,
31'b0011110000000000000010000000000,
31'b1100000000001000000000000100100,
31'b0100000010000010000000010000010,
31'b0100000010000000000000010000010,
31'b0010000000000001000000100100000,
31'b1100000000000000000000000100100,
31'b0100000000100000000001100000000,
31'b0000001000000001000000000001000,
31'b1000001010000000000000000010001,
31'b1000000100000000000000001000100,
31'b0100000000011000000001100000000,
31'b1010000001000000100000000000001,
31'b0000101000010000000000000000100,
31'b1000000100001000000000001000100,
31'b0100000000010000000001100000000,
31'b0100000000100000000110000010000,
31'b0000101000001000000000000000100,
31'b1000000100010000000000001000100,
31'b0100000000001000000001100000000,
31'b0100000010100000000000010000010,
31'b0000101000000000000000000000100,
31'b1000000000000000000000100001001,
31'b0100000000000000000001100000000,
31'b0100000000000010000001100000000,
31'b0000100000000100000000001100010,
31'b0000100000000000010000110000000,
31'b0000100000000000000000001100010,
31'b0100000001010000000000010000010,
31'b0101001000100000000001000000000,
31'b0001000000000001000000100001000,
31'b0011001000000001000000000100000,
31'b0011000000000000000001000000101,
31'b0000000000000011001000000100000,
31'b0000000000000001001000000100000,
31'b0100100000000000001000100000001,
31'b0100000001000000000000010000010,
31'b1010000000000000000100001100000,
31'b1000010000000000000000010001000,
31'b1000010100000000010100000000000,
31'b1000010000000100000000010001000,
31'b1110000100000000000100000000000,
31'b0010000110000000011000000000000,
31'b0001100000001000000000100000100,
31'b1100001000000000000000001000010,
31'b0101001000000000000001000000000,
31'b0101001000000010000001000000000,
31'b0001100000000000000000100000100,
31'b1001001000000000000000000001001,
31'b1010000000000000001000000001001,
31'b0010000000000000100100010000000,
31'b0110000000000010001001000000000,
31'b0110000000000000001001000000000,
31'b0101001000010000000001000000000,
31'b1000010000100000000000010001000,
31'b0100100100000000000000000000010,
31'b0110000000001000001001000000000,
31'b0000000000000101000000100010000,
31'b0100100000000000000000000110001,
31'b0000000000000001000000100010000,
31'b0100000000010000000000010000010,
31'b0000001000000001101000000000000,
31'b0001000100000000100001001000000,
31'b0000001000100000000010000000010,
31'b0100000010000000000110000010000,
31'b0100000000000110000000010000010,
31'b0100000000000100000000010000010,
31'b0100000000000010000000010000010,
31'b0100000000000000000000010000010,
31'b0010100100000000100100000000000,
31'b1100000010000000000000000100100,
31'b0100000010100000000001100000000,
31'b0100000000001000000000010000010,
31'b1000001000000000000000000010001,
31'b1000001000000010000000000010001,
31'b0000001000001000000010000000010,
31'b0100001000000000000001000011000,
31'b0000000100000000010000100000000,
31'b0000011000000000000000001001000,
31'b0000001000000000000010000000010,
31'b0000001000000010000010000000010,
31'b1000110100000000000000000001000,
31'b0101000000000000100001000100000,
31'b0100000010001000000001100000000,
31'b0100000000100000000000010000010,
31'b0000101010000000000000000000100,
31'b1000010000000000010000000010100,
31'b0100000010000000000001100000000,
31'b0100000010000010000001100000000,
31'b0111100000000000000000000000000,
31'b0111100000000010000000000000000,
31'b1100000100000000001000001000000,
31'b0000010010000000000010010000010,
31'b0111100000001000000000000000000,
31'b1000010000000000000010000100100,
31'b1000000100000000000100100000100,
31'b0000010000010000000100000010000,
31'b0111100000010000000000000000000,
31'b0100000000000000000101001000000,
31'b1000000000101000001000000100000,
31'b0000010000001000000100000010000,
31'b1000000001000000000111000000000,
31'b0000010000000100000100000010000,
31'b1000000000100000001000000100000,
31'b0000010000000000000100000010000,
31'b1010000010000000001000000010000,
31'b1011001000000000000000000100000,
31'b1001000000000000000000100001000,
31'b1001000000000010000000100001000,
31'b1000000001000010000000100010000,
31'b1000000001000000000000100010000,
31'b1000000000010000001000000100000,
31'b1000000001000100000000100010000,
31'b1000001011000000000000000001000,
31'b0100100000000000010010000000001,
31'b1000000000001000001000000100000,
31'b1010000000000000100000000011000,
31'b1000000000000100001000000100000,
31'b1000000001010000000000100010000,
31'b1000000000000000001000000100000,
31'b1000000000000010001000000100000,
31'b0111100001000000000000000000000,
31'b1000001000000001000010000000010,
31'b0110000100000000010000000000100,
31'b0000000100001000001010000000000,
31'b1000000000100010000000100010000,
31'b1000000000100000000000100010000,
31'b0000000100000010001010000000000,
31'b0000000100000000001010000000000,
31'b0010000010000000000001000000100,
31'b0100100010000000000000000101000,
31'b0011000000000000010000100000010,
31'b0001010100000000010000010000000,
31'b1000000000000000000111000000000,
31'b1000000000110000000000100010000,
31'b1000000001100000001000000100000,
31'b0000010001000000000100000010000,
31'b1000001010010000000000000001000,
31'b1000000000001000000000100010000,
31'b1001000001000000000000100001000,
31'b1000001000000000101000000000000,
31'b1000000000000010000000100010000,
31'b1000000000000000000000100010000,
31'b1000000001010000001000000100000,
31'b1000000000000100000000100010000,
31'b1000001010000000000000000001000,
31'b1000001010000010000000000001000,
31'b1000001010000100000000000001000,
31'b1010000010000000000000100100000,
31'b0000010100000000000000000000100,
31'b1000000000010000000000100010000,
31'b1000000001000000001000000100000,
31'b1000000001000010001000000100000,
31'b0000000000000000000000011001000,
31'b0010010000000000000100000100000,
31'b0010000100000000000010100000000,
31'b0000010000000000000010010000010,
31'b0010000000000001100000000000001,
31'b1000010000000000000000010010001,
31'b0010000100001000000010100000000,
31'b0001000001000000000000011010000,
31'b0010000001000000000001000000100,
31'b0100100001000000000000000101000,
31'b0010000100010000000010100000000,
31'b0001000100000000100010000010000,
31'b0010000001001000000001000000100,
31'b0010010000000000000000000000111,
31'b1000101000000000010100000000000,
31'b0001000000000000011000000000010,
31'b1010000000000000001000000010000,
31'b1010000000000010001000000010000,
31'b1010000000000100001000000010000,
31'b0100010000000001000101000000000,
31'b1010000000001000001000000010000,
31'b1000000000000000100000000101000,
31'b1010001000000000100000100000000,
31'b1001001000010000000000000010000,
31'b1000001001000000000000000001000,
31'b1001000000000000101000100000000,
31'b1000001001000100000000000001000,
31'b1010000001000000000000100100000,
31'b1000001001001000000000000001000,
31'b1001001000000100000000000010000,
31'b1000000010000000001000000100000,
31'b1001001000000000000000000010000,
31'b0010000000010000000001000000100,
31'b0101010000000000000001010000000,
31'b0010000101000000000010100000000,
31'b0001010000000000101100000000000,
31'b0010000001000001100000000000001,
31'b1100000000000000000010010001000,
31'b0000000100000001000000001000100,
31'b0001000000000000000000011010000,
31'b0010000000000000000001000000100,
31'b0100100000000000000000000101000,
31'b0010000000000100000001000000100,
31'b1010000000100000000000100100000,
31'b0010000000001000000001000000100,
31'b0100100000001000000000000101000,
31'b0010000000001100000001000000100,
31'b0001000001000000011000000000010,
31'b1000001000010000000000000001000,
31'b1000001000010010000000000001000,
31'b1001000000000000100000000110000,
31'b1010000000010000000000100100000,
31'b1000001000011000000000000001000,
31'b1000000010000000000000100010000,
31'b0100010000000000010001000000100,
31'b1011000000000000001000000001000,
31'b1000001000000000000000000001000,
31'b1000001000000010000000000001000,
31'b1000001000000100000000000001000,
31'b1010000000000000000000100100000,
31'b1000001000001000000000000001000,
31'b1000001000001010000000000001000,
31'b1000001000001100000000000001000,
31'b1010000000001000000000100100000,
31'b1100000000000100001000001000000,
31'b0000001010000000000010000101000,
31'b1100000000000000001000001000000,
31'b0000000010000000010100001000000,
31'b1000010000000000001001000010000,
31'b0000000001000100001010000000000,
31'b1000000000000000000100100000100,
31'b0000000001000000001010000000000,
31'b0011001001000000000010000000000,
31'b1100100000000001000000000000010,
31'b1100000000010000001000001000000,
31'b0001010001000000010000010000000,
31'b0000010001100000000000000000100,
31'b0000010100000100000100000010000,
31'b1000000100100000001000000100000,
31'b0000010100000000000100000010000,
31'b0000010001011000000000000000100,
31'b0000001001000000010000000000001,
31'b1100000000100000001000001000000,
31'b0000101000000000001000001100000,
31'b0000010001010000000000000000100,
31'b0000000000000000000101000100000,
31'b1000000100010000001000000100000,
31'b0000000001100000001010000000000,
31'b0000010001001000000000000000100,
31'b0000010000000001010100000000000,
31'b1100000000000000000000000001110,
31'b0010000010000000000101000010000,
31'b0000010001000000000000000000100,
31'b0000010001000010000000000000100,
31'b1000000100000000001000000100000,
31'b1000000100000010001000000100000,
31'b0110000000000100010000000000100,
31'b0000001000100000010000000000001,
31'b0110000000000000010000000000100,
31'b0000000000001000001010000000000,
31'b0000010000110000000000000000100,
31'b0000000000000100001010000000000,
31'b0000000000000010001010000000000,
31'b0000000000000000001010000000000,
31'b0011001000000000000010000000000,
31'b0011001000000010000010000000000,
31'b0110000000010000010000000000100,
31'b0001010000000000010000010000000,
31'b0000010000100000000000000000100,
31'b0000010000100010000000000000100,
31'b0000010000100100000000000000100,
31'b0000000000010000001010000000000,
31'b0000010000011000000000000000100,
31'b0000001000000000010000000000001,
31'b0110000000100000010000000000100,
31'b0000001000000100010000000000001,
31'b0000010000010000000000000000100,
31'b0000000000000001100000000000010,
31'b0000010000010100000000000000100,
31'b0000000000100000001010000000000,
31'b0000010000001000000000000000100,
31'b0000010000001010000000000000100,
31'b0100001000000000001000010000000,
31'b0101000000000000000010000000101,
31'b0000010000000000000000000000100,
31'b0000010000000010000000000000100,
31'b0000010000000100000000000000100,
31'b0000010000000110000000000000100,
31'b0010000000000100000010100000000,
31'b0000001000000000000010000101000,
31'b0010000000000000000010100000000,
31'b0000000000000000010100001000000,
31'b0010000100000001100000000000001,
31'b0000101000000000011001000000000,
31'b0010000000001000000010100000000,
31'b0000000011000000001010000000000,
31'b0010000101000000000001000000100,
31'b1100000000000000100000001001000,
31'b0010000000010000000010100000000,
31'b0001000000000000100010000010000,
31'b0000000001000000100010000001000,
31'b1001000000000000100000000000011,
31'b0010000000011000000010100000000,
31'b0001000100000000011000000000010,
31'b1100100000000000000010000001000,
31'b0000100001001000000000001001000,
31'b0010000000100000000010100000000,
31'b0000100000000000000011000000001,
31'b0101110000000000000001000000000,
31'b0000100001000000000000001001000,
31'b0010001000000001000000000010010,
31'b0000100001000100000000001001000,
31'b1100010000000001001000000000000,
31'b0010010000000000001000100000100,
31'b0010000000110000000010100000000,
31'b0010000000000000000101000010000,
31'b0100000000000000000000010101000,
31'b0110010000000000000100001000000,
31'b1000001000000001000000010000100,
31'b1001001100000000000000000010000,
31'b0010000100010000000001000000100,
31'b0000100000101000000000001001000,
31'b0010000001000000000010100000000,
31'b0000000010001000001010000000000,
31'b0000000000010000100010000001000,
31'b0000100000100000000000001001000,
31'b0000000000000001000000001000100,
31'b0000000010000000001010000000000,
31'b0010000100000000000001000000100,
31'b0100100100000000000000000101000,
31'b0010000100000100000001000000100,
31'b0001010010000000010000010000000,
31'b0000000000000000100010000001000,
31'b0000100000000000001000000000110,
31'b0000000000010001000000001000100,
31'b0000010000000000100000001000010,
31'b1000110000000000000000000010001,
31'b0000100000001000000000001001000,
31'b0010010000000000000000000110100,
31'b0000100001000000000011000000001,
31'b0000100000000010000000001001000,
31'b0000100000000000000000001001000,
31'b0000110000000000000010000000010,
31'b0000100000000100000000001001000,
31'b1000001100000000000000000001000,
31'b1000010000000000010000101000000,
31'b1000010000000000000000010100010,
31'b1010000100000000000000100100000,
31'b0000010010000000000000000000100,
31'b0000100000010000000000001001000,
31'b0000010010000100000000000000100,
31'b0000100000010100000000001001000,
31'b0010000010000000010000000000010,
31'b1011000000100000000000000100000,
31'b0011000000000000000001100000100,
31'b1101000000000001000001000000000,
31'b0100000000000001000000001000010,
31'b0100100000010100001000000000000,
31'b0100100000010010001000000000000,
31'b0100100000010000001000000000000,
31'b1000000011100000000000000001000,
31'b0100100000001100001000000000000,
31'b0110000100000000000001000000010,
31'b0100100000001000001000000000000,
31'b0100100000000110001000000000000,
31'b0100100000000100001000000000000,
31'b0100100000000010001000000000000,
31'b0100100000000000001000000000000,
31'b1011000000000010000000000100000,
31'b1011000000000000000000000100000,
31'b1001001000000000000000100001000,
31'b1000000001000000101000000000000,
31'b0100110000000000000010000000100,
31'b1011000000001000000000000100000,
31'b1010000010000000100000100000000,
31'b1001000010010000000000000010000,
31'b1000000011000000000000000001000,
31'b1011000000010000000000000100000,
31'b1000001000001000001000000100000,
31'b1001000010001000000000000010000,
31'b1000001000000100001000000100000,
31'b1010000000000000001000100001000,
31'b1000001000000000001000000100000,
31'b1001000010000000000000000010000,
31'b1000000010110000000000000001000,
31'b1000000000000001000010000000010,
31'b1000010000000001000000001001000,
31'b1000000000100000101000000000000,
31'b0100100000000000000000100110000,
31'b0000000000000101000000000010001,
31'b0000000000000011000000000010001,
31'b0000000000000001000000000010001,
31'b1000000010100000000000000001000,
31'b1000000010100010000000000001000,
31'b1000100000000000001010001000000,
31'b1000100010000001000000000000100,
31'b1000001000000000000111000000000,
31'b0100100001000100001000000000000,
31'b0100100001000010001000000000000,
31'b0100100001000000001000000000000,
31'b1000000010010000000000000001000,
31'b0000000100000000010000000000001,
31'b1000000000000010101000000000000,
31'b1000000000000000101000000000000,
31'b1000001000000010000000100010000,
31'b1000001000000000000000100010000,
31'b1010000000000000000000000111000,
31'b1000000000001000101000000000000,
31'b1000000010000000000000000001000,
31'b1000000010000010000000000001000,
31'b1000000010000100000000000001000,
31'b1000000000010000101000000000000,
31'b1000000010001000000000000001000,
31'b1000001000010000000000100010000,
31'b1000001001000000001000000100000,
31'b1001000011000000000000000010000,
31'b0010000000000000010000000000010,
31'b0010000000000010010000000000010,
31'b0010000000000100010000000000010,
31'b0010000000000110010000000000010,
31'b0100100000000000100000000001000,
31'b0100100000000010100000000001000,
31'b1010000000100000100000100000000,
31'b1001000000110000000000000010000,
31'b1000000001100000000000000001000,
31'b1001000100000001010000000000000,
31'b1000100000001000010100000000000,
31'b1001000000101000000000000010000,
31'b1000100000000100010100000000000,
31'b1001000000100100000000000010000,
31'b1000100000000000010100000000000,
31'b1001000000100000000000000010000,
31'b1000000001010000000000000001000,
31'b1011000010000000000000000100000,
31'b1010000000001000100000100000000,
31'b1001000000011000000000000010000,
31'b1010000000000100100000100000000,
31'b1001000000010100000000000010000,
31'b1010000000000000100000100000000,
31'b1001000000010000000000000010000,
31'b1000000001000000000000000001000,
31'b1000000001000010000000000001000,
31'b1000000001000100000000000001000,
31'b1001000000001000000000000010000,
31'b1000000001001000000000000001000,
31'b1001000000000100000000000010000,
31'b0100010000000000000000000000010,
31'b1001000000000000000000000010000,
31'b1000000000110000000000000001000,
31'b1000000010000001000010000000010,
31'b1000110000000000100000000000010,
31'b1000100000010001000000000000100,
31'b1100000000000000000100100000010,
31'b0010010000000000010001000000001,
31'b0001000100000000000010000110000,
31'b0001000000000000001001000000100,
31'b1000000000100000000000000001000,
31'b1000000000100010000000000001000,
31'b1000000000100100000000000001000,
31'b1000100000000001000000000000100,
31'b1000000000101000000000000001000,
31'b1000000000101010000000000001000,
31'b1000100001000000010100000000000,
31'b1001000001100000000000000010000,
31'b1000000000010000000000000001000,
31'b1000000000010010000000000001000,
31'b1000000000010100000000000001000,
31'b1000000010000000101000000000000,
31'b1000000000011000000000000001000,
31'b1000001010000000000000100010000,
31'b1010000001000000100000100000000,
31'b1001000001010000000000000010000,
31'b1000000000000000000000000001000,
31'b1000000000000010000000000001000,
31'b1000000000000100000000000001000,
31'b0100000000000000000001000000001,
31'b1000000000001000000000000001000,
31'b1000000000001010000000000001000,
31'b1000000000001100000000000001000,
31'b1001000001000000000000000010000,
31'b0011000001010000000010000000000,
31'b0000000010000000000010000101000,
31'b1100001000000000001000001000000,
31'b0000100000100000001000001100000,
31'b1100100000000000000101000000000,
31'b0000100010000000011001000000000,
31'b1000100000000000101000010000000,
31'b0000100000000000000100000001001,
31'b0011000001000000000010000000000,
31'b1010000000000000000000000001011,
31'b0110000000000000000001000000010,
31'b0110000000000010000001000000010,
31'b0011000001001000000010000000000,
31'b1111000000000000000000001000000,
31'b0110000000001000000001000000010,
31'b0100100100000000001000000000000,
31'b0000000001000010010000000000001,
31'b0000000001000000010000000000001,
31'b0100000001010000001000010000000,
31'b0000100000000000001000001100000,
31'b0000010000000000010001000000010,
31'b0000001000000000000101000100000,
31'b0010000010000001000000000010010,
31'b0000100000100000000100000001001,
31'b0000000000000001000000000100010,
31'b0000000001010000010000000000001,
31'b0100000001000000001000010000000,
31'b0100100000000000000000100000011,
31'b0000011001000000000000000000100,
31'b0000011001000010000000000000100,
31'b1000001100000000001000000100000,
31'b1001000110000000000000000010000,
31'b0011000000010000000010000000000,
31'b0000000000100000010000000000001,
31'b0110001000000000010000000000100,
31'b0000001000001000001010000000000,
31'b0011000000011000000010000000000,
31'b0000001000000100001010000000000,
31'b0001000000000000000000010000101,
31'b0000001000000000001010000000000,
31'b0011000000000000000010000000000,
31'b0011000000000010000010000000000,
31'b0100000000100000001000010000000,
31'b0110010000001000000000000000001,
31'b0011000000001000000010000000000,
31'b0110010000000100000000000000001,
31'b0110010000000010000000000000001,
31'b0110010000000000000000000000001,
31'b0000000000000010010000000000001,
31'b0000000000000000010000000000001,
31'b0100000000010000001000010000000,
31'b0000000000000100010000000000001,
31'b0000011000010000000000000000100,
31'b0000000000001000010000000000001,
31'b0101010000000000010010000000000,
31'b0000001000100000001010000000000,
31'b0000000000000000100101000000000,
31'b0000000000010000010000000000001,
31'b0100000000000000001000010000000,
31'b0100000000000010001000010000000,
31'b0000011000000000000000000000100,
31'b0000011000000010000000000000100,
31'b0100000000001000001000010000000,
31'b0110010000100000000000000000001,
31'b0010000100000000010000000000010,
31'b0000000000000000000010000101000,
31'b0010001000000000000010100000000,
31'b0000001000000000010100001000000,
31'b0100100100000000100000000001000,
31'b0000100000000000011001000000000,
31'b0010001000001000000010100000000,
31'b0000100010000000000100000001001,
31'b1001000000000011010000000000000,
31'b1001000000000001010000000000000,
31'b0110000010000000000001000000010,
31'b1001000000000101010000000000000,
31'b1001000001000000000100000000100,
31'b1000100000000000000000010001000,
31'b1000100100000000010100000000000,
31'b1001000100100000000000000010000,
31'b1010000000000001000010000000001,
31'b0000000011000000010000000000001,
31'b0010001000100000000010100000000,
31'b0000101000000000000011000000001,
31'b0010000000000101000000000010010,
31'b0000101001000000000000001001000,
31'b0010000000000001000000000010010,
31'b1001000100010000000000000010000,
31'b1000000101000000000000000001000,
31'b1001000000100001010000000000000,
31'b1000000101000100000000000001000,
31'b1001000100001000000000000010000,
31'b1000000101001000000000000001000,
31'b1001000100000100000000000010000,
31'b1000000000000001000000010000100,
31'b1001000100000000000000000010000,
31'b1001000000000000000000000100011,
31'b0000000010100000010000000000001,
31'b0011100000000000000000000000110,
31'b0000001010001000001010000000000,
31'b1100000000000000000000001101000,
31'b0000101000100000000000001001000,
31'b0001000000000000000010000110000,
31'b0000001010000000001010000000000,
31'b1000000100100000000000000001000,
31'b1001000001000001010000000000000,
31'b1001100000000000000000010010000,
31'b1000100100000001000000000000100,
31'b1001000000000000000100000000100,
31'b1001000000000010000100000000100,
31'b1001000000000100000100000000100,
31'b0110010010000000000000000000001,
31'b1000000100010000000000000001000,
31'b0000000010000000010000000000001,
31'b1000000100010100000000000001000,
31'b0000000010000100010000000000001,
31'b1000000100011000000000000001000,
31'b0000101000000000000000001001000,
31'b0010100000000000000000101100000,
31'b0000101000000100000000001001000,
31'b1000000100000000000000000001000,
31'b1000000100000010000000000001000,
31'b1000000100000100000000000001000,
31'b1000000000000000010100010000000,
31'b1000000100001000000000000001000,
31'b1000100000000000010000000010100,
31'b1000000100001100000000000001000,
31'b1001000101000000000000000010000,
31'b0111110000000000000000000000000,
31'b0010000010000000000100000100000,
31'b0000001010000000000100100001000,
31'b0000000010000000000010010000010,
31'b1000000100000000001001000010000,
31'b1000000000000000000010000100100,
31'b0000000000100000000011100000000,
31'b0000000000010000000100000010000,
31'b0001000001000000000100000001000,
31'b0000100000000000000000010000100,
31'b0000000000100001000000010001000,
31'b0000000000001000000100000010000,
31'b0000000101100000000000000000100,
31'b0000000000000100000100000010000,
31'b0000000000000010000100000010000,
31'b0000000000000000000100000010000,
31'b0000000101011000000000000000100,
31'b0010101000000000011000000000000,
31'b0000000000010001000000010001000,
31'b0100000010000001000101000000000,
31'b0000000101010000000000000000100,
31'b1000010001000000000000100010000,
31'b0000000000000000000011100000000,
31'b0000000000110000000100000010000,
31'b0000000101001000000000000000100,
31'b0000100000100000000000010000100,
31'b0000000000000001000000010001000,
31'b0000000000101000000100000010000,
31'b0000000101000000000000000000100,
31'b0000000101000010000000000000100,
31'b0001100000000000010000000000000,
31'b0000000000100000000100000010000,
31'b0100000000000000000000001100100,
31'b0101000010000000000001010000000,
31'b1101000000000000110000000000000,
31'b0001000100010000010000010000000,
31'b0000000100110000000000000000100,
31'b1000010000100000000000100010000,
31'b0000010100000010001010000000000,
31'b0000010100000000001010000000000,
31'b0001000000000000000100000001000,
31'b0001000000000010000100000001000,
31'b0001000000000100000100000001000,
31'b0001000100000000010000010000000,
31'b0000000100100000000000000000100,
31'b0000000100100010000000000000100,
31'b0000000100100100000000000000100,
31'b0000000001000000000100000010000,
31'b0000000100011000000000000000100,
31'b1000101000000000000000001000100,
31'b0010000100000000000010010000001,
31'b1100000000000000000001101000000,
31'b0000000100010000000000000000100,
31'b1000010000000000000000100010000,
31'b0000000100010100000000000000100,
31'b1000010000000100000000100010000,
31'b0000000100001000000000000000100,
31'b0000100000000000010000000011000,
31'b0000000100001100000000000000100,
31'b0001100000000001000100000000100,
31'b0000000100000000000000000000100,
31'b0000000100000010000000000000100,
31'b0000000100000100000000000000100,
31'b0000000100000110000000000000100,
31'b0010000000000010000100000100000,
31'b0010000000000000000100000100000,
31'b0000001000000000000100100001000,
31'b0000000000000000000010010000010,
31'b1000000000000010000000010010001,
31'b1000000000000000000000010010001,
31'b0100001000110000000000000000010,
31'b0000000010010000000100000010000,
31'b0010010001000000000001000000100,
31'b0010000000010000000100000100000,
31'b0100001000101000000000000000010,
31'b0000000010001000000100000010000,
31'b0100001000100100000000000000010,
31'b0010000000000000000000000000111,
31'b0100001000100000000000000000010,
31'b0000000010000000000100000010000,
31'b1010010000000000001000000010000,
31'b0010000000100000000100000100000,
31'b0100001000011000000000000000010,
31'b0100000000000001000101000000000,
31'b0101100100000000000001000000000,
31'b1000010000000000100000000101000,
31'b0100001000010000000000000000010,
31'b0100001000010010000000000000010,
31'b1100000100000001001000000000000,
31'b0010000100000000001000100000100,
31'b0100001000001000000000000000010,
31'b0100001000001010000000000000010,
31'b0100001000000100000000000000010,
31'b0110000100000000000100001000000,
31'b0100001000000000000000000000010,
31'b0100001000000010000000000000010,
31'b0101000000000010000001010000000,
31'b0101000000000000000001010000000,
31'b1001000000000000000000010001001,
31'b0001000000000000101100000000000,
31'b0010001000010000100100000000000,
31'b1100000000000000010000100100000,
31'b1100000000000000000000011000010,
31'b0001010000000000000000011010000,
31'b0010010000000000000001000000100,
31'b0101000000010000000001010000000,
31'b0010010000000100000001000000100,
31'b0001000110000000010000010000000,
31'b0010001000000000100100000000000,
31'b0010001000000010100100000000000,
31'b0110000000000000000000001010100,
31'b0000000100000000100000001000010,
31'b1000100100000000000000000010001,
31'b0101000000100000000001010000000,
31'b0100000000001000010001000000100,
31'b0100000000000000100000000100010,
31'b0000101000000000010000100000000,
31'b1000010010000000000000100010000,
31'b0100000000000000010001000000100,
31'b0100000000001000100000000100010,
31'b1000011000000000000000000001000,
31'b1000011000000010000000000001000,
31'b1000011000000100000000000001000,
31'b1010010000000000000000100100000,
31'b0000000110000000000000000000100,
31'b0000001000000000000000001010001,
31'b0100001001000000000000000000010,
31'b0100001001000010000000000000010,
31'b1100100000000000100000000000100,
31'b0010100000000001100000100000000,
31'b1100010000000000001000001000000,
31'b0001000001010000010000010000000,
31'b1000000000000000001001000010000,
31'b1000000100000000000010000100100,
31'b1000010000000000000100100000100,
31'b0000010001000000001010000000000,
31'b0001100000000001000000000010000,
31'b0000100100000000000000010000100,
31'b0001100000000101000000000010000,
31'b0001000001000000010000010000000,
31'b0000000001100000000000000000100,
31'b0000000100000100000100000010000,
31'b0000000100000010000100000010000,
31'b0000000100000000000100000010000,
31'b0000000001011000000000000000100,
31'b0000001000000000100000000100100,
31'b0010000001000000000010010000001,
31'b1100000000000001100000000001000,
31'b0000000001010000000000000000100,
31'b0000010000000000000101000100000,
31'b0000000100000000000011100000000,
31'b0000010001100000001010000000000,
31'b0000000001001000000000000000100,
31'b0000000000000001010100000000000,
31'b0000000100000001000000010001000,
31'b0001000000000000000000000011100,
31'b0000000001000000000000000000100,
31'b0000000001000010000000000000100,
31'b0000000001000100000000000000100,
31'b0000000100100000000100000010000,
31'b0101000000000000001000000000001,
31'b0101000000000010001000000000001,
31'b0110010000000000010000000000100,
31'b0001000000010000010000010000000,
31'b0000000000110000000000000000100,
31'b0000010000000100001010000000000,
31'b0000010000000010001010000000000,
31'b0000010000000000001010000000000,
31'b0000000000101000000000000000100,
31'b0001000000000100010000010000000,
31'b0001000000000010010000010000000,
31'b0001000000000000010000010000000,
31'b0000000000100000000000000000100,
31'b0000000000100010000000000000100,
31'b0000000000100100000000000000100,
31'b0000100000000001000000000001000,
31'b0000000000011000000000000000100,
31'b0000011000000000010000000000001,
31'b0010000000000000000010010000001,
31'b0011001000000000001000000000100,
31'b0000000000010000000000000000100,
31'b0000000000010010000000000000100,
31'b0000000000010100000000000000100,
31'b0000010000100000001010000000000,
31'b0000000000001000000000000000100,
31'b0000000000001010000000000000100,
31'b0000000000001100000000000000100,
31'b0001000000100000010000010000000,
31'b0000000000000000000000000000100,
31'b0000000000000010000000000000100,
31'b0000000000000100000000000000100,
31'b0000000000000110000000000000100,
31'b0010010000000100000010100000000,
31'b0010000100000000000100000100000,
31'b0010010000000000000010100000000,
31'b0000010000000000010100001000000,
31'b1001000000000001000000000000101,
31'b1001001000000000000001000100000,
31'b0011100000000001000000000100000,
31'b0000010011000000001010000000000,
31'b1100000000100001001000000000000,
31'b0010000100010000000100000100000,
31'b1100000000000000100010000000010,
31'b0001010000000000100010000010000,
31'b0100000000000000100000000010001,
31'b0110000000100000000100001000000,
31'b0100001100100000000000000000010,
31'b0000000110000000000100000010000,
31'b1100000000010001001000000000000,
31'b0010000100100000000100000100000,
31'b0010010000100000000010100000000,
31'b1100100000000000000000001000010,
31'b0101100000000000000001000000000,
31'b0110000000010000000100001000000,
31'b0001001000000000000000100000100,
31'b1001100000000000000000000001001,
31'b1100000000000001001000000000000,
31'b0010000000000000001000100000100,
31'b1100000000000101001000000000000,
31'b0010010000000000000101000010000,
31'b0000000011000000000000000000100,
31'b0110000000000000000100001000000,
31'b0100001100000000000000000000010,
31'b0110000000000100000100001000000,
31'b1001000000010000100001000000000,
31'b1010000000000000000001100010000,
31'b0010010001000000000010100000000,
31'b0001000100000000101100000000000,
31'b0000100000000001101000000000000,
31'b0000110000100000000000001001000,
31'b0000100000100000000010000000010,
31'b0000010010000000001010000000000,
31'b1001000000000000100001000000000,
31'b1001000000000010100001000000000,
31'b1001000000000100100001000000000,
31'b0001000010000000010000010000000,
31'b0000000010100000000000000000100,
31'b0000000010100010000000000000100,
31'b0000000010100100000000000000100,
31'b0000000000000000100000001000010,
31'b1000100000000000000000000010001,
31'b1000100000000010000000000010001,
31'b0010000000000000000000000110100,
31'b0100100000000000000001000011000,
31'b0000000010010000000000000000100,
31'b0000110000000000000000001001000,
31'b0000100000000000000010000000010,
31'b0000100000000010000010000000010,
31'b0000000010001000000000000000100,
31'b1000000000000000010000101000000,
31'b1000000000000000000000010100010,
31'b1000000000000100010000101000000,
31'b0000000010000000000000000000100,
31'b0000000010000010000000000000100,
31'b0000000010000100000000000000100,
31'b0000000010000110000000000000100,
31'b0011000000000000001100000010000,
31'b0010100000100000011000000000000,
31'b0000000010000000000100100001000,
31'b0100000000010000000001110000000,
31'b1000000100000000000000011000100,
31'b1001000000000001000000001010000,
31'b0100000010110000000000000000010,
31'b0100000000000001000010000001000,
31'b1000000001000000100010000000100,
31'b0000101000000000000000010000100,
31'b0100000010101000000000000000010,
31'b0100000000000000000001110000000,
31'b0100000010100100000000000000010,
31'b0100000000000000100000001000100,
31'b0100000010100000000000000000010,
31'b0000001000000000000100000010000,
31'b0110000000000000000000000110010,
31'b0010100000000000011000000000000,
31'b0100000010011000000000000000010,
31'b1001000100000000010000001000000,
31'b0100100000000000000010000000100,
31'b0100100000000010000010000000100,
31'b0100000010010000000000000000010,
31'b0100000010010010000000000000010,
31'b1100000000000000000000010100100,
31'b0010100000010000011000000000000,
31'b0100000010001000000000000000010,
31'b0100000010001010000000000000010,
31'b0100000010000100000000000000010,
31'b0100000010000110000000000000010,
31'b0100000010000000000000000000010,
31'b0100000010000010000000000000010,
31'b1000000000010000100010000000100,
31'b1000100000100000000000001000100,
31'b1000000000000001000000001001000,
31'b1000010000100000101000000000000,
31'b0010000100000000011000010000000,
31'b0010000010000000010001000000001,
31'b1010000000000000100000010000001,
31'b0010000000000000001100000001000,
31'b1000000000000000100010000000100,
31'b1000100000000000001000000001010,
31'b1000000000010001000000001001000,
31'b0110000100001000000000000000001,
31'b0010000010000000100100000000000,
31'b0110000100000100000000000000001,
31'b0110000100000010000000000000001,
31'b0110000100000000000000000000001,
31'b1000100000000010000000001000100,
31'b1000100000000000000000001000100,
31'b1000010000000010101000000000000,
31'b1000010000000000101000000000000,
31'b0000100010000000010000100000000,
31'b1000100000001000000000001000100,
31'b0101000100000000010010000000000,
31'b1000010000001000101000000000000,
31'b1000010010000000000000000001000,
31'b1000100000010000000000001000100,
31'b1000010010000100000000000001000,
31'b1000010000010000101000000000000,
31'b0000001100000000000000000000100,
31'b0000001100000010000000000000100,
31'b0100000011000000000000000000010,
31'b0110000100100000000000000000001,
31'b0010010000000000010000000000010,
31'b0010001000000000000100000100000,
31'b0000000000000000000100100001000,
31'b0000001000000000000010010000010,
31'b0100110000000000100000000001000,
31'b1001000100000000000001000100000,
31'b0100000000110000000000000000010,
31'b0100000010000001000010000001000,
31'b1100000000000000110000100000000,
31'b0010001000010000000100000100000,
31'b0100000000101000000000000000010,
31'b0100000010000000000001110000000,
31'b0100000000100100000000000000010,
31'b0100000010000000100000001000100,
31'b0100000000100000000000000000010,
31'b0100000000100010000000000000010,
31'b1110100000000000000100000000000,
31'b0010100010000000011000000000000,
31'b0100000000011000000000000000010,
31'b0100001000000001000101000000000,
31'b0100000000010100000000000000010,
31'b0100100000000001001000001000000,
31'b0100000000010000000000000000010,
31'b0100000000010010000000000000010,
31'b1000010001000000000000000001000,
31'b1101000000000000000001001000000,
31'b0100000000001000000000000000010,
31'b0100000000001010000000000000010,
31'b0100000000000100000000000000010,
31'b0100000000000110000000000000010,
31'b0100000000000000000000000000010,
31'b0100000000000010000000000000010,
31'b1000100000000100100000000000010,
31'b0101001000000000000001010000000,
31'b1000100000000000100000000000010,
31'b1000100000000010100000000000010,
31'b0010000000010000100100000000000,
31'b0010000000000000010001000000001,
31'b1110000000000000010000000001000,
31'b0010000010000000001100000001000,
31'b1000010000100000000000000001000,
31'b1000010000100010000000000001000,
31'b1000100000010000100000000000010,
31'b1000110000000001000000000000100,
31'b0010000000000000100100000000000,
31'b0010000000000010100100000000000,
31'b0100000001100000000000000000010,
31'b0110000110000000000000000000001,
31'b1000010000010000000000000001000,
31'b1000100010000000000000001000100,
31'b1000100000100000100000000000010,
31'b1000010010000000101000000000000,
31'b0000100000000000010000100000000,
31'b0000100000000010010000100000000,
31'b0100000001010000000000000000010,
31'b0100000001010010000000000000010,
31'b1000010000000000000000000001000,
31'b1000010000000010000000000001000,
31'b1000010000000100000000000001000,
31'b1000000000000000000010001000010,
31'b0001000000000000000011000000000,
31'b0000000000000000000000001010001,
31'b0100000001000000000000000000010,
31'b0100000001000010000000000000010,
31'b1000000000001000000000011000100,
31'b0000000010000000010000110000000,
31'b1000000000000000100001100000000,
31'b1001000000100000010000001000000,
31'b1000000000000000000000011000100,
31'b1001000010000000000001000100000,
31'b1000000000001000100001100000000,
31'b0110000001010000000000000000001,
31'b0011010001000000000010000000000,
31'b0000101100000000000000010000100,
31'b1010000000000000000010001000001,
31'b1011000000000000000001000010000,
31'b0010000000000000000000001010010,
31'b0110000001000100000000000000001,
31'b0110000001000010000000000000001,
31'b0110000001000000000000000000001,
31'b0000000000001000010001000000010,
31'b0000000000000000100000000100100,
31'b1001000000000010010000001000000,
31'b1001000000000000010000001000000,
31'b0000000000000000010001000000010,
31'b0000000000001000100000000100100,
31'b0001000010000000000000100000100,
31'b1001000000001000010000001000000,
31'b0000010000000001000000000100010,
31'b0000001000000001010100000000000,
31'b0100010001000000001000010000000,
31'b1001000000010000010000001000000,
31'b0000001001000000000000000000100,
31'b0000001001000010000000000000100,
31'b0100000110000000000000000000010,
31'b0110000001100000000000000000001,
31'b0101001000000000001000000000001,
31'b0100000000000000000010010000100,
31'b1000000100000001000000001001000,
31'b0110000000011000000000000000001,
31'b0010000000000000011000010000000,
31'b0110000000010100000000000000001,
31'b0110000000010010000000000000001,
31'b0110000000010000000000000000001,
31'b0011010000000000000010000000000,
31'b0110000000001100000000000000001,
31'b0110000000001010000000000000001,
31'b0110000000001000000000000000001,
31'b0000001000100000000000000000100,
31'b0110000000000100000000000000001,
31'b0110000000000010000000000000001,
31'b0110000000000000000000000000001,
31'b0000010000000010010000000000001,
31'b0000010000000000010000000000001,
31'b0101000000001000010010000000000,
31'b0011000000000000001000000000100,
31'b0000001000010000000000000000100,
31'b0000010000001000010000000000001,
31'b0101000000000000010010000000000,
31'b0110000000110000000000000000001,
31'b0000001000001000000000000000100,
31'b0000010000010000010000000000001,
31'b0100010000000000001000010000000,
31'b0110000000101000000000000000001,
31'b0000001000000000000000000000100,
31'b0000001000000010000000000000100,
31'b0000001000000100000000000000100,
31'b0110000000100000000000000000001,
31'b0000000000000100000000001100010,
31'b0000000000000000010000110000000,
31'b0000000000000000000000001100010,
31'b0000000000000100010000110000000,
31'b1001000000000010000001000100000,
31'b1001000000000000000001000100000,
31'b0001000000100000000000100000100,
31'b1001000000000100000001000100000,
31'b0100000000000100001000100000001,
31'b0000100000000001001000000100000,
31'b0100000000000000001000100000001,
31'b0100100001000000000000010000010,
31'b0100001000000000100000000010001,
31'b1001000000010000000001000100000,
31'b0100000100100000000000000000010,
31'b0110000011000000000000000000001,
31'b0001000000001100000000100000100,
31'b0000000010000000100000000100100,
31'b0001000000001000000000100000100,
31'b1001000010000000010000001000000,
31'b0001000000000100000000100000100,
31'b1001000000100000000001000100000,
31'b0001000000000000000000100000100,
31'b1000000000000000100000010000010,
31'b1100001000000001001000000000000,
31'b0010100000000000100100010000000,
31'b0100000100001000000000000000010,
31'b0110100000000000001001000000000,
31'b0100000100000100000000000000010,
31'b0110001000000000000100001000000,
31'b0100000100000000000000000000010,
31'b0100000100000010000000000000010,
31'b0100000000000010000000000110001,
31'b0100000000000000000000000110001,
31'b0000100000000001000000100010000,
31'b0100100000010000000000010000010,
31'b0010000100010000100100000000000,
31'b1110000000000000000100010000000,
31'b0001010000000000000010000110000,
31'b1100000000000000000010000100010,
31'b1001001000000000100001000000000,
31'b0100100000000100000000010000010,
31'b0100100000000010000000010000010,
31'b0100100000000000000000010000010,
31'b0010000100000000100100000000000,
31'b0110000010000100000000000000001,
31'b0110000010000010000000000000001,
31'b0110000010000000000000000000001,
31'b1000101000000000000000000010001,
31'b0000010010000000010000000000001,
31'b0011000000000001000010001000000,
31'b0011000010000000001000000000100,
31'b0000100100000000010000100000000,
31'b0000111000000000000000001001000,
31'b0001000001000000000000100000100,
31'b1001000000000000001110000000000,
31'b1000010100000000000000000001000,
31'b1000010100000010000000000001000,
31'b1000010100000100000000000001000,
31'b1000010000000000010100010000000,
31'b0000001010000000000000000000100,
31'b0000001010000010000000000000100,
31'b0100000101000000000000000000010,
31'b0110000010100000000000000000001,
31'b1000000000000000000000000000000,
31'b1000000000000010000000000000000,
31'b1000000000000100000000000000000,
31'b1000000000000110000000000000000,
31'b1000000000001000000000000000000,
31'b1000000000001010000000000000000,
31'b1000000000001100000000000000000,
31'b1000000000001110000000000000000,
31'b1000000000010000000000000000000,
31'b1000000000010010000000000000000,
31'b1000000000010100000000000000000,
31'b1000000000010110000000000000000,
31'b1000000000011000000000000000000,
31'b1000000000011010000000000000000,
31'b1000000000011100000000000000000,
31'b1011001000000000001000000000000,
31'b1000000000100000000000000000000,
31'b1000000000100010000000000000000,
31'b1000000000100100000000000000000,
31'b1000000000100110000000000000000,
31'b1000000000101000000000000000000,
31'b1000000000101010000000000000000,
31'b1000000000101100000000000000000,
31'b1001000000000000010000010000100,
31'b1000000000110000000000000000000,
31'b1000000000110010000000000000000,
31'b1000000000110100000000000000000,
31'b1000010000000000001010000000100,
31'b1000000000111000000000000000000,
31'b1100001000000000000010010000000,
31'b1110010000000000010000000000000,
31'b0011000000000000010000000010010,
31'b1000000001000000000000000000000,
31'b1000000001000010000000000000000,
31'b1000000001000100000000000000000,
31'b1000000001000110000000000000000,
31'b1000000001001000000000000000000,
31'b0100000000000000000010001000000,
31'b1000000001001100000000000000000,
31'b1001000000000000000000000011000,
31'b1000000001010000000000000000000,
31'b1000000001010010000000000000000,
31'b1000000001010100000000000000000,
31'b1000000001010110000000000000000,
31'b1000000001011000000000000000000,
31'b1000001000000000100000000100000,
31'b1010000000000000100000100001000,
31'b1001000000010000000000000011000,
31'b1000000001100000000000000000000,
31'b1000000001100010000000000000000,
31'b1000000001100100000000000000000,
31'b1000000100000000000100000010100,
31'b1000000001101000000000000000000,
31'b1000100100000000000000010000000,
31'b1000100000000000010100000001000,
31'b1001000000100000000000000011000,
31'b0000001000000000000000011000000,
31'b0000000100000000000010000100000,
31'b0000010000000000000100100000000,
31'b0000010000000010000100100000000,
31'b0100100000000000100000000000000,
31'b0100100000000010100000000000000,
31'b0100100000000100100000000000000,
31'b0100100000000110100000000000000,
31'b1000000010000000000000000000000,
31'b1000000010000010000000000000000,
31'b1000000010000100000000000000000,
31'b1000000010000110000000000000000,
31'b1000000010001000000000000000000,
31'b1000000010001010000000000000000,
31'b1000000010001100000000000000000,
31'b1001000000000000100000100100000,
31'b1000000010010000000000000000000,
31'b1000000010010010000000000000000,
31'b0000000000000000000100010000001,
31'b1000000000000000101000000001000,
31'b1000000010011000000000000000000,
31'b1000001000000000000000100011000,
31'b1010000000000000000000000110000,
31'b1010000000000010000000000110000,
31'b1000000010100000000000000000000,
31'b1000000010100010000000000000000,
31'b1000000010100100000000000000000,
31'b1000000010100110000000000000000,
31'b1000000010101000000000000000000,
31'b1000000010101010000000000000000,
31'b1000000010101100000000000000000,
31'b0100100001000000001000000001000,
31'b1000000010110000000000000000000,
31'b1000000010110010000000000000000,
31'b1000010000000001000000001000000,
31'b1000010000000011000000001000000,
31'b1100000000000001000001000010000,
31'b0010010000000100001100000000000,
31'b1010000000100000000000000110000,
31'b0010010000000000001100000000000,
31'b1000000011000000000000000000000,
31'b1000000011000010000000000000000,
31'b1000000011000100000000000000000,
31'b1010001000000000100000000010000,
31'b1000000011001000000000000000000,
31'b1010000000000000001000100000000,
31'b1000001000000000001000000101000,
31'b1010000000000100001000100000000,
31'b1000000011010000000000000000000,
31'b1011000000000000000000000101000,
31'b1001001000000000000000100000000,
31'b1001001000000010000000100000000,
31'b1001000000000000101000000010000,
31'b1010000000010000001000100000000,
31'b1010000001000000000000000110000,
31'b0100100000000000000000001000110,
31'b1000000011100000000000000000000,
31'b1010000100000000000000000000011,
31'b1000001000000000000100001000001,
31'b0100100000001000001000000001000,
31'b1000100000000000001001000000001,
31'b1010000000100000001000100000000,
31'b0100100000000010001000000001000,
31'b0100100000000000001000000001000,
31'b0001000000000001000000000000001,
31'b0001000000000011000000000000001,
31'b0001000000000101000000000000001,
31'b0101100000000000000000100100000,
31'b0100100010000000100000000000000,
31'b0100100010000010100000000000000,
31'b0100100010000100100000000000000,
31'b0100010000000001000010000000000,
31'b1000000100000000000000000000000,
31'b1000000100000010000000000000000,
31'b1000000100000100000000000000000,
31'b1000000100000110000000000000000,
31'b1000000100001000000000000000000,
31'b1000000100001010000000000000000,
31'b1000000100001100000000000000000,
31'b1001100000000001000100000000000,
31'b1000000100010000000000000000000,
31'b0100000000000000100000010000000,
31'b1000000100010100000000000000000,
31'b0000000000000000001101000000000,
31'b1000000100011000000000000000000,
31'b0000101000000000000000001000000,
31'b1010000000000001000001001000000,
31'b0000101000000100000000001000000,
31'b1000000100100000000000000000000,
31'b1000000100100010000000000000000,
31'b1000000100100100000000000000000,
31'b1000000100100110000000000000000,
31'b0000001000000000100010000000000,
31'b1000100001000000000000010000000,
31'b1000000000000001010000000010000,
31'b1000100001000100000000010000000,
31'b1000000100110000000000000000000,
31'b0000000001000000000010000100000,
31'b1000010000000000000001000110000,
31'b0000000001000100000010000100000,
31'b1100000000000000000000001100000,
31'b0000101000100000000000001000000,
31'b1100000000000100000000001100000,
31'b0000101000100100000000001000000,
31'b1000000101000000000000000000000,
31'b1000000101000010000000000000000,
31'b1000000101000100000000000000000,
31'b1000000101000110000000000000000,
31'b1000000101001000000000000000000,
31'b1000100000100000000000010000000,
31'b1000000101001100000000000000000,
31'b1001000100000000000000000011000,
31'b1000000101010000000000000000000,
31'b0000000000100000000010000100000,
31'b1000000101010100000000000000000,
31'b0000000001000000001101000000000,
31'b1000000101011000000000000000000,
31'b0000101001000000000000001000000,
31'b0010000010000000000101100000000,
31'b0000101001000100000000001000000,
31'b1000000101100000000000000000000,
31'b0000000000010000000010000100000,
31'b1000000101100100000000000000000,
31'b1000000000000000000100000010100,
31'b1000100000000010000000010000000,
31'b1000100000000000000000010000000,
31'b1000100000000110000000010000000,
31'b1000100000000100000000010000000,
31'b0000000000000010000010000100000,
31'b0000000000000000000010000100000,
31'b0000010100000000000100100000000,
31'b0000000000000100000010000100000,
31'b0100100100000000100000000000000,
31'b0000000000001000000010000100000,
31'b0101010000000000000000000100001,
31'b0000100010000000000100000000001,
31'b1000000110000000000000000000000,
31'b1000000110000010000000000000000,
31'b1000000110000100000000000000000,
31'b1100000000000000100100000000001,
31'b1000000110001000000000000000000,
31'b1000110000000000000000100000001,
31'b1100010000000001000000000100000,
31'b0010010000000000000000100100100,
31'b1000000110010000000000000000000,
31'b0000000000000000010000000001001,
31'b1100000000000000010001000000000,
31'b0000000010000000001101000000000,
31'b1000010000000000010000001010000,
31'b0000101010000000000000001000000,
31'b1100000000001000010001000000000,
31'b0000101010000100000000001000000,
31'b1000000110100000000000000000000,
31'b1010000001000000000000000000011,
31'b1110000000000000000000001010000,
31'b0011010000000000000000001000010,
31'b1010010000000000000001000000000,
31'b1010010000000010000001000000000,
31'b1010010000000100000001000000000,
31'b0010000001000000000010000010000,
31'b1010000000000001010000000100000,
31'b0000000011000000000010000100000,
31'b1100000000100000010001000000000,
31'b0000101000000000010001000100000,
31'b1100000010000000000000001100000,
31'b0000101010100000000000001000000,
31'b0001000001000000100010100000000,
31'b0000100001000000000100000000001,
31'b1000000111000000000000000000000,
31'b1010000000100000000000000000011,
31'b1100001000000000000000000000110,
31'b0010001000000001000000100000010,
31'b1000010000000000001000010000010,
31'b1010000100000000001000100000000,
31'b0010000000100010000010000010000,
31'b0010000000100000000010000010000,
31'b1001000000000000010010000000010,
31'b0000000010100000000010000100000,
31'b1100000001000000010001000000000,
31'b0000100000101000000100000000001,
31'b0010010000000000001000000010100,
31'b0000101011000000000000001000000,
31'b0010000000000000000101100000000,
31'b0000100000100000000100000000001,
31'b1010000000000010000000000000011,
31'b1010000000000000000000000000011,
31'b0110000000000000000001000001010,
31'b0010000000001000000010000010000,
31'b1010010001000000000001000000000,
31'b1000100010000000000000010000000,
31'b0010000000000010000010000010000,
31'b0010000000000000000010000010000,
31'b0001000100000001000000000000001,
31'b0000000010000000000010000100000,
31'b0001000100000101000000000000001,
31'b0000100000001000000100000000001,
31'b0100100110000000100000000000000,
31'b0000100000000100000100000000001,
31'b0001000000000000100010100000000,
31'b0000100000000000000100000000001,
31'b1000001000000000000000000000000,
31'b1000001000000010000000000000000,
31'b1000001000000100000000000000000,
31'b1000001000000110000000000000000,
31'b1000001000001000000000000000000,
31'b1000001000001010000000000000000,
31'b1000001000001100000000000000000,
31'b1011000000010000001000000000000,
31'b1000001000010000000000000000000,
31'b1000001000010010000000000000000,
31'b1000001000010100000000000000000,
31'b1011000000001000001000000000000,
31'b1000001000011000000000000000000,
31'b0000100100000000000000001000000,
31'b1011000000000010001000000000000,
31'b1011000000000000001000000000000,
31'b1000001000100000000000000000000,
31'b0100100000000000000000000100000,
31'b0000000000000001000000100000001,
31'b0100100000000100000000000100000,
31'b0000000100000000100010000000000,
31'b0100100000001000000000000100000,
31'b0000000100000100100010000000000,
31'b0100100000001100000000000100000,
31'b0000000001000000000000011000000,
31'b0100100000010000000000000100000,
31'b0000000001000100000000011000000,
31'b0100100000010100000000000100000,
31'b0000000100010000100010000000000,
31'b1100000000000000000010010000000,
31'b0000000100010100100010000000000,
31'b1100000000000100000010010000000,
31'b1000001001000000000000000000000,
31'b1000001001000010000000000000000,
31'b1000001001000100000000000000000,
31'b1010000010000000100000000010000,
31'b1000001001001000000000000000000,
31'b1000000000010000100000000100000,
31'b1000001001001100000000000000000,
31'b1001001000000000000000000011000,
31'b0000000000100000000000011000000,
31'b1000000000001000100000000100000,
31'b1001000010000000000000100000000,
31'b1001000010000010000000100000000,
31'b1000000000000010100000000100000,
31'b1000000000000000100000000100000,
31'b1001000010001000000000100000000,
31'b1000000000000100100000000100000,
31'b0000000000010000000000011000000,
31'b0100100001000000000000000100000,
31'b0000000001000001000000100000001,
31'b0100100001000100000000000100000,
31'b0000000101000000100010000000000,
31'b1000101100000000000000010000000,
31'b0010000100000001000001010000000,
31'b0011000000000000000001000010100,
31'b0000000000000000000000011000000,
31'b0000000000000010000000011000000,
31'b0000000000000100000000011000000,
31'b0000000000000110000000011000000,
31'b0000000000001000000000011000000,
31'b1000000000100000100000000100000,
31'b0000000000001100000000011000000,
31'b1001000000000000000001010000010,
31'b1000001010000000000000000000000,
31'b1000001010000010000000000000000,
31'b1000001010000100000000000000000,
31'b1010000001000000100000000010000,
31'b1000001010001000000000000000000,
31'b1000001010001010000000000000000,
31'b1000001010001100000000000000000,
31'b0100100000000000010001001000000,
31'b1000001010010000000000000000000,
31'b1000001010010010000000000000000,
31'b1001000001000000000000100000000,
31'b1001000001000010000000100000000,
31'b1000001010011000000000000000000,
31'b1000000000000000000000100011000,
31'b1010001000000000000000000110000,
31'b1011000010000000001000000000000,
31'b0001010000000000000100000000000,
31'b0100100010000000000000000100000,
31'b0001010000000100000100000000000,
31'b0100100010000100000000000100000,
31'b0001010000001000000100000000000,
31'b0100100010001000000000000100000,
31'b0101100000000000100000100000000,
31'b0100000000000000000110000000001,
31'b0001010000010000000100000000000,
31'b0110000000000000000100010000100,
31'b1001000001100000000000100000000,
31'b0110100000001000000000000010000,
31'b0001010000011000000100000000000,
31'b1100000010000000000010010000000,
31'b0110100000000010000000000010000,
31'b0110100000000000000000000010000,
31'b1000001011000000000000000000000,
31'b1010000000000100100000000010000,
31'b0000010000000001000000010000000,
31'b1010000000000000100000000010000,
31'b1000001011001000000000000000000,
31'b1010001000000000001000100000000,
31'b1000000000000000001000000101000,
31'b1010000000001000100000000010000,
31'b1001000000000100000000100000000,
31'b1001000000000110000000100000000,
31'b1001000000000000000000100000000,
31'b1001000000000010000000100000000,
31'b1001000000001100000000100000000,
31'b1000000010000000100000000100000,
31'b1001000000001000000000100000000,
31'b1001000000001010000000100000000,
31'b0001010001000000000100000000000,
31'b0100100011000000000000000100000,
31'b1000000000000000000100001000001,
31'b1010000000100000100000000010000,
31'b0001010001001000000100000000000,
31'b0010000000000101001000000000001,
31'b1000000000100000001000000101000,
31'b0010000000000001001000000000001,
31'b0000000010000000000000011000000,
31'b0001000000000000000001000100100,
31'b1001000000100000000000100000000,
31'b1001000000100010000000100000000,
31'b0001000000000000110000000000010,
31'b1000000010100000100000000100000,
31'b1001000000101000000000100000000,
31'b0110100001000000000000000010000,
31'b1000001100000000000000000000000,
31'b1000001100000010000000000000000,
31'b1000001100000100000000000000000,
31'b1010000000000000000100001000010,
31'b0000000000100000100010000000000,
31'b0000100000010000000000001000000,
31'b0000000000000001001000000000010,
31'b0000100000010100000000001000000,
31'b1000001100010000000000000000000,
31'b0000100000001000000000001000000,
31'b1001100000000000000001000000010,
31'b0000100000001100000000001000000,
31'b0000100000000010000000001000000,
31'b0000100000000000000000001000000,
31'b0000100000000110000000001000000,
31'b0000100000000100000000001000000,
31'b0000000000001000100010000000000,
31'b0100100100000000000000000100000,
31'b0000000100000001000000100000001,
31'b0101010000000000100000000000001,
31'b0000000000000000100010000000000,
31'b0000000000000010100010000000000,
31'b0000000000000100100010000000000,
31'b0000110010000001000000000000000,
31'b0000000101000000000000011000000,
31'b0000100000101000000000001000000,
31'b0010000001000000000010100001000,
31'b0000100010000000010001000100000,
31'b0000000000010000100010000000000,
31'b0000100000100000000000001000000,
31'b0000000000010100100010000000000,
31'b0000100000100100000000001000000,
31'b1000001101000000000000000000000,
31'b1100000000100000100000001000000,
31'b1100000010000000000000000000110,
31'b0010000010000001000000100000010,
31'b0100000000000000000000010100000,
31'b0100000000000010000000010100000,
31'b0100000000000100000000010100000,
31'b0100000000000110000000010100000,
31'b1100100000000000000010000000000,
31'b0000100001001000000000001000000,
31'b1100100000000100000010000000000,
31'b0000100001001100000000001000000,
31'b0100000000010000000000010100000,
31'b0000100001000000000000001000000,
31'b0100100000000000000000000010011,
31'b0000100001000100000000001000000,
31'b0000000100010000000000011000000,
31'b1100000000000000100000001000000,
31'b0010000000010000000010100001000,
31'b1100000000000100100000001000000,
31'b0000000001000000100010000000000,
31'b1000101000000000000000010000000,
31'b0010000000000001000001010000000,
31'b1000101000000100000000010000000,
31'b0000000100000000000000011000000,
31'b0000001000000000000010000100000,
31'b0010000000000000000010100001000,
31'b0000001000000100000010000100000,
31'b0000000100001000000000011000000,
31'b0000100001100000000000001000000,
31'b0010000000010001000001010000000,
31'b0000101010000000000100000000001,
31'b1000001110000000000000000000000,
31'b1000001110000010000000000000000,
31'b1100000001000000000000000000110,
31'b0010100000000000000000001110000,
31'b0000010000000000000000000001100,
31'b0000100010010000000000001000000,
31'b0000010000000100000000000001100,
31'b0000110000100001000000000000000,
31'b1000100000000000010000100000100,
31'b0000100010001000000000001000000,
31'b1100001000000000010001000000000,
31'b0000100010001100000000001000000,
31'b0000100010000010000000001000000,
31'b0000100010000000000000001000000,
31'b0000100010000110000000001000000,
31'b0000100010000100000000001000000,
31'b0001010100000000000100000000000,
31'b0100100110000000000000000100000,
31'b0001010100000100000100000000000,
31'b0001000000000000000010100100000,
31'b0000000010000000100010000000000,
31'b0000110000000101000000000000000,
31'b0000110000000011000000000000000,
31'b0000110000000001000000000000000,
31'b0001010100010000000100000000000,
31'b0000100010101000000000001000000,
31'b0110000000000000010000000001100,
31'b0000100000000000010001000100000,
31'b0000010000000000001000001000010,
31'b0000100010100000000000001000000,
31'b0000100000000000100000000000110,
31'b0000000000000000001010000001000,
31'b1100000000000100000000000000110,
31'b0010000000000101000000100000010,
31'b1100000000000000000000000000110,
31'b0010000000000001000000100000010,
31'b0100000010000000000000010100000,
31'b0101000000000000000001001000100,
31'b1100000000001000000000000000110,
31'b0010001000100000000010000010000,
31'b1100100010000000000010000000000,
31'b0000100011001000000000001000000,
31'b1001000100000000000000100000000,
31'b1100010000000001100000000000000,
31'b0110100000000000000100000000100,
31'b0000100011000000000000001000000,
31'b1100000000000000000100000100001,
31'b0000101000100000000100000000001,
31'b0001010101000000000100000000000,
31'b1100000010000000100000001000000,
31'b1100000000100000000000000000110,
31'b0010001000001000000010000010000,
31'b0000010000000000010000010010000,
31'b1010000000000001110000000000000,
31'b0010001000000010000010000010000,
31'b0010001000000000000010000010000,
31'b0001000000000000001010000010000,
31'b0000001010000000000010000100000,
31'b1100000000000000001000001001000,
31'b0000101000001000000100000000001,
31'b0001000100000000110000000000010,
31'b0000101000000100000100000000001,
31'b1001000000000000001000000000011,
31'b0000101000000000000100000000001,
31'b1000010000000000000000000000000,
31'b1000010000000010000000000000000,
31'b1000010000000100000000000000000,
31'b1000010000000110000000000000000,
31'b1000010000001000000000000000000,
31'b1000010000001010000000000000000,
31'b1000010000001100000000000000000,
31'b1101000000000000000010000000001,
31'b1000010000010000000000000000000,
31'b1000010000010010000000000000000,
31'b1000010000010100000000000000000,
31'b1000010000010110000000000000000,
31'b1000010000011000000000000000000,
31'b1000010000011010000000000000000,
31'b1110000000100000010000000000000,
31'b0010101000000000010000000100000,
31'b1000010000100000000000000000000,
31'b1000010000100010000000000000000,
31'b1000010000100100000000000000000,
31'b1000010000100110000000000000000,
31'b1000010000101000000000000000000,
31'b1010000000000000001000010000001,
31'b1110000000010000010000000000000,
31'b0010000100000000110000010000000,
31'b1000010000110000000000000000000,
31'b1000010000110010000000000000000,
31'b0000000001000000000100100000000,
31'b1000000000000000001010000000100,
31'b1110000000000100010000000000000,
31'b0010000010000100001100000000000,
31'b1110000000000000010000000000000,
31'b0010000010000000001100000000000,
31'b1000010001000000000000000000000,
31'b1000010001000010000000000000000,
31'b0001000000000000000000001000001,
31'b0000000000000000000011000010000,
31'b1000010001001000000000000000000,
31'b1000000000000000000001000000011,
31'b0100000000000000000000000001010,
31'b0100000000000010000000000001010,
31'b1000010001010000000000000000000,
31'b1000010001010010000000000000000,
31'b0000000000100000000100100000000,
31'b0000000000100010000100100000000,
31'b1000010001011000000000000000000,
31'b1000011000000000100000000100000,
31'b0100000000010000000000000001010,
31'b0100000010100001000010000000000,
31'b1000010001100000000000000000000,
31'b1000010001100010000000000000000,
31'b0000000000010000000100100000000,
31'b0000000000100000000011000010000,
31'b1010100000000000000000100000010,
31'b1000110100000000000000010000000,
31'b0100000000100000000000000001010,
31'b0100000010010001000010000000000,
31'b0000000000000100000100100000000,
31'b0000010100000000000010000100000,
31'b0000000000000000000100100000000,
31'b0000000000000010000100100000000,
31'b0100110000000000100000000000000,
31'b0100110000000010100000000000000,
31'b0000000000001000000100100000000,
31'b0100000010000001000010000000000,
31'b1000010010000000000000000000000,
31'b1000010010000010000000000000000,
31'b1000010010000100000000000000000,
31'b1000100000000001100010000000000,
31'b1000010010001000000000000000000,
31'b1000100100000000000000100000001,
31'b1100000100000001000000000100000,
31'b0010000100000000000000100100100,
31'b1000010010010000000000000000000,
31'b1000100000000000000000001001100,
31'b1000000000100001000000001000000,
31'b1000010000000000101000000001000,
31'b1000010010011000000000000000000,
31'b0101000000000000000110010000000,
31'b1010010000000000000000000110000,
31'b0010000000100000001100000000000,
31'b0001001000000000000100000000000,
31'b1000100000000000001000000000010,
31'b1000000000010001000000001000000,
31'b1000100000000100001000000000010,
31'b1010000100000000000001000000000,
31'b1010000100000010000001000000000,
31'b1010000100000100000001000000000,
31'b0010000000010000001100000000000,
31'b1000000000000101000000001000000,
31'b1000100000010000001000000000010,
31'b1000000000000001000000001000000,
31'b1000000000000011000000001000000,
31'b1010000100010000000001000000000,
31'b0010000000000100001100000000000,
31'b1000000000001001000000001000000,
31'b0010000000000000001100000000000,
31'b1000010011000000000000000000000,
31'b1010100000000000000001010000000,
31'b0000001000000001000000010000000,
31'b0000001000000011000000010000000,
31'b1000010011001000000000000000000,
31'b1010010000000000001000100000000,
31'b0100000010000000000000000001010,
31'b0100000010000010000000000001010,
31'b1001000000000000000100011000000,
31'b0100000100000000010010000010000,
31'b0000001000010001000000010000000,
31'b0100001000000000000000100010010,
31'b0100100000000000000010000001100,
31'b0100000000000000101000000000010,
31'b0100000010010000000000000001010,
31'b0100000000100001000010000000000,
31'b1000000000000000000000110000001,
31'b1000100001000000001000000000010,
31'b0000001000100001000000010000000,
31'b0100000000011001000010000000000,
31'b1010000101000000000001000000000,
31'b0100000000010101000010000000000,
31'b0100000010100000000000000001010,
31'b0100000000010001000010000000000,
31'b0001010000000001000000000000001,
31'b0100000100000000100000100000001,
31'b0000000010000000000100100000000,
31'b0100000000001001000010000000000,
31'b0100110010000000100000000000000,
31'b0100000000000101000010000000000,
31'b0100000000000011000010000000000,
31'b0100000000000001000010000000000,
31'b1000010100000000000000000000000,
31'b1000010100000010000000000000000,
31'b1000010100000100000000000000000,
31'b1000010100000110000000000000000,
31'b1000010100001000000000000000000,
31'b1000100010000000000000100000001,
31'b1100000010000001000000000100000,
31'b0010000010000000000000100100100,
31'b1000010100010000000000000000000,
31'b0000000000000000000000100010100,
31'b1000010100010100000000000000000,
31'b0000010000000000001101000000000,
31'b1000010100011000000000000000000,
31'b0000111000000000000000001000000,
31'b0001000001000000000000100001100,
31'b0000100000000000000100110000000,
31'b1000010100100000000000000000000,
31'b1000010100100010000000000000000,
31'b1000010100100100000000000000000,
31'b0101001000000000100000000000001,
31'b1010000010000000000001000000000,
31'b1010000010000010000001000000000,
31'b1010000010000100000001000000000,
31'b0010000000000000110000010000000,
31'b1000010100110000000000000000000,
31'b0000010001000000000010000100000,
31'b1000000000000000000001000110000,
31'b1000000100000000001010000000100,
31'b1100010000000000000000001100000,
31'b0001100001000001000000100000000,
31'b1110000100000000010000000000000,
31'b0010000110000000001100000000000,
31'b1000010101000000000000000000000,
31'b1000010101000010000000000000000,
31'b0000000000000000001000000100100,
31'b0000000100000000000011000010000,
31'b1000010101001000000000000000000,
31'b1000110000100000000000010000000,
31'b0100000100000000000000000001010,
31'b0110000000000000010010000100000,
31'b1000010101010000000000000000000,
31'b0000010000100000000010000100000,
31'b0000000100100000000100100000000,
31'b0000010001000000001101000000000,
31'b0011000000000001000001000000001,
31'b0011001000000000000000000100100,
31'b0001000000000000000000100001100,
31'b1001101000000000000000000000001,
31'b1000010101100000000000000000000,
31'b1000000000000000001001100000000,
31'b0000000100010000000100100000000,
31'b1000010000000000000100000010100,
31'b1010000011000000000001000000000,
31'b1000110000000000000000010000000,
31'b0101000000010000000000000100001,
31'b1000110000000100000000010000000,
31'b0000010000000010000010000100000,
31'b0000010000000000000010000100000,
31'b0000000100000000000100100000000,
31'b0000010000000100000010000100000,
31'b0101000000000100000000000100001,
31'b0001100000000001000000100000000,
31'b0101000000000000000000000100001,
31'b0101000000000010000000000100001,
31'b1000010110000000000000000000000,
31'b1000100000001000000000100000001,
31'b1100000000001001000000000100000,
31'b0011000000100000000000001000010,
31'b0000001000000000000000000001100,
31'b1000100000000000000000100000001,
31'b1100000000000001000000000100000,
31'b0010000000000000000000100100100,
31'b1000010110010000000000000000000,
31'b0000010000000000010000000001001,
31'b1100010000000000010001000000000,
31'b0011000000000000001000000001100,
31'b1000000000000000010000001010000,
31'b1000100000010000000000100000001,
31'b1100000000010001000000000100000,
31'b0010000100100000001100000000000,
31'b1010000000001000000001000000000,
31'b1010000000001010000001000000000,
31'b1010000000001100000001000000000,
31'b0011000000000000000000001000010,
31'b1010000000000000000001000000000,
31'b1010000000000010000001000000000,
31'b1010000000000100000001000000000,
31'b0000101000000001000000000000000,
31'b1010000000011000000001000000000,
31'b0100000001000000100000100000001,
31'b1000000100000001000000001000000,
31'b1001001000000000001001000000000,
31'b1010000000010000000001000000000,
31'b1010000000010010000001000000000,
31'b1010000000010100000001000000000,
31'b0010000100000000001100000000000,
31'b1000010111000000000000000000000,
31'b0101000000000000100100001000000,
31'b0000001100000001000000010000000,
31'b0001001000000000000000000010100,
31'b1000000000000000001000010000010,
31'b1000100001000000000000100000001,
31'b1100000001000001000000000100000,
31'b0010010000100000000010000010000,
31'b0110100000000000100001000000000,
31'b0100000000000000010010000010000,
31'b0010100000000000001100010000000,
31'b1100001000000001100000000000000,
31'b0010000000000000001000000010100,
31'b0100000100000000101000000000010,
31'b0010010000000000000101100000000,
31'b1100000000000000010000000000011,
31'b1010000001001000000001000000000,
31'b1010010000000000000000000000011,
31'b0000101000000000010100000000100,
31'b0011000001000000000000001000010,
31'b1010000001000000000001000000000,
31'b1010000001000010000001000000000,
31'b1010000001000100000001000000000,
31'b0010010000000000000010000010000,
31'b0101100000000000000110000000000,
31'b0100000000000000100000100000001,
31'b0000100000000001100000000100000,
31'b0100000100001001000010000000000,
31'b1010000001010000000001000000000,
31'b0100000100000101000010000000000,
31'b0101000010000000000000000100001,
31'b0100000100000001000010000000000,
31'b1000011000000000000000000000000,
31'b1000011000000010000000000000000,
31'b1000011000000100000000000000000,
31'b1010000000000000010010010000000,
31'b1000011000001000000000000000000,
31'b1000011000001010000000000000000,
31'b1100000000000000001000010000100,
31'b0010100000010000010000000100000,
31'b1000011000010000000000000000000,
31'b1000011000010010000000000000000,
31'b1001000000100000000000010000001,
31'b0100100100000000000001000010000,
31'b1000011000011000000000000000000,
31'b1000000000000000010000000000101,
31'b0110000000000000001000000010010,
31'b0010100000000000010000000100000,
31'b0001000010000000000100000000000,
31'b0100110000000000000000000100000,
31'b0001000010000100000100000000000,
31'b0101000100000000100000000000001,
31'b0001000010001000000100000000000,
31'b0101000000000001000010100000000,
31'b0001100000000000000010000100001,
31'b0000100110000001000000000000000,
31'b0001000010010000000100000000000,
31'b0101000000000000000001010001000,
31'b1001000000000000000000010000001,
31'b1001000000000010000000010000001,
31'b0001000010011000000100000000000,
31'b1100010000000000000010010000000,
31'b1110001000000000010000000000000,
31'b0010100000100000010000000100000,
31'b1000011001000000000000000000000,
31'b1000011001000010000000000000000,
31'b0000000010000001000000010000000,
31'b0000001000000000000011000010000,
31'b1000011001001000000000000000000,
31'b1000010000010000100000000100000,
31'b0100001000000000000000000001010,
31'b0100001000000010000000000001010,
31'b1000000000000001000100000000001,
31'b1000010000001000100000000100000,
31'b0000001000100000000100100000000,
31'b0100000010000000000000100010010,
31'b1000010000000010100000000100000,
31'b1000010000000000100000000100000,
31'b0100001000010000000000000001010,
31'b1001100100000000000000000000001,
31'b0001000011000000000100000000000,
31'b0111000000000000000000001000100,
31'b0000001000010000000100100000000,
31'b0000001000100000000011000010000,
31'b0001000011001000000100000000000,
31'b0011000000000000001100100000000,
31'b0100001000100000000000000001010,
31'b0000000010000000000100000011000,
31'b0000010000000000000000011000000,
31'b0010000000000000000100000101000,
31'b0000001000000000000100100000000,
31'b0000001000000010000100100000000,
31'b0000010000001000000000011000000,
31'b1000010000100000100000000100000,
31'b0100000000000000000001010010000,
31'b0100001010000001000010000000000,
31'b0001000000100000000100000000000,
31'b0000100000000000010000000010000,
31'b0000000001000001000000010000000,
31'b0000100000000100010000000010000,
31'b0000000100000000000000000001100,
31'b0000100000001000010000000010000,
31'b0000000100000100000000000001100,
31'b0000100100100001000000000000000,
31'b0000000000000000000000101000001,
31'b0000100000010000010000000010000,
31'b0000000001010001000000010000000,
31'b0100100000000001000000001100000,
31'b0000000100010000000000000001100,
31'b1000010000000000000000100011000,
31'b0000000100010100000000000001100,
31'b0010100010000000010000000100000,
31'b0001000000000000000100000000000,
31'b0001000000000010000100000000000,
31'b0001000000000100000100000000000,
31'b0001000000000110000100000000000,
31'b0001000000001000000100000000000,
31'b0001000000001010000100000000000,
31'b0001000000001100000100000000000,
31'b0000100100000001000000000000000,
31'b0001000000010000000100000000000,
31'b0010100000000000000001001000000,
31'b1000001000000001000000001000000,
31'b1001000100000000001001000000000,
31'b0001000000011000000100000000000,
31'b0010100000001000000001001000000,
31'b1011100000000000000000000000010,
31'b0010001000000000001100000000000,
31'b0000000000000101000000010000000,
31'b0000100001000000010000000010000,
31'b0000000000000001000000010000000,
31'b0000000000000011000000010000000,
31'b0000000101000000000000000001100,
31'b0001100100000000000100010000000,
31'b0000000000001001000000010000000,
31'b0000000000100000000100000011000,
31'b0000000001000000000000101000001,
31'b0100000000000100000000100010010,
31'b0000000000010001000000010000000,
31'b0100000000000000000000100010010,
31'b0010000100000000000001011000000,
31'b1100000000000000000010100000001,
31'b0000000000011001000000010000000,
31'b0100001000100001000010000000000,
31'b0001000001000000000100000000000,
31'b0001000001000010000100000000000,
31'b0000000000100001000000010000000,
31'b0000000000100011000000010000000,
31'b0001000001001000000100000000000,
31'b0001000000000001010000000000100,
31'b0000000000101001000000010000000,
31'b0000000000000000000100000011000,
31'b0001000001010000000100000000000,
31'b0010100001000000000001001000000,
31'b0000001010000000000100100000000,
31'b0100001000001001000010000000000,
31'b0001010000000000110000000000010,
31'b1100000000000000110000000010000,
31'b0100001000000011000010000000000,
31'b0100001000000001000010000000000,
31'b1000011100000000000000000000000,
31'b1000011100000010000000000000000,
31'b1000011100000100000000000000000,
31'b0101000000100000100000000000001,
31'b0000000010000000000000000001100,
31'b0000110000010000000000001000000,
31'b0000010000000001001000000000010,
31'b0000100010100001000000000000000,
31'b1000100000000000000000000011001,
31'b0000110000001000000000001000000,
31'b0110000000000000110010000000000,
31'b0100100000000000000001000010000,
31'b0000110000000010000000001000000,
31'b0000110000000000000000001000000,
31'b0000100000000000000010000001010,
31'b0000000000000000101000000000100,
31'b0001000110000000000100000000000,
31'b0101000000000100100000000000001,
31'b0101000000000010100000000000001,
31'b0101000000000000100000000000001,
31'b0000010000000000100010000000000,
31'b0000100010000101000000000000000,
31'b0000100010000011000000000000000,
31'b0000100010000001000000000000000,
31'b0001000110010000000100000000000,
31'b0010100000000001000000000110000,
31'b1001000100000000000000010000001,
31'b1001000010000000001001000000000,
31'b0000010000010000100010000000000,
31'b0000110000100000000000001000000,
31'b0000100010010011000000000000000,
31'b0000100010010001000000000000000,
31'b1100000000000001001000000001000,
31'b0011000000000000000100000000011,
31'b0000001000000000001000000100100,
31'b0001000010000000000000000010100,
31'b0100010000000000000000010100000,
31'b0110000000000000000100001001000,
31'b0100010000000100000000010100000,
31'b1001100000010000000000000000001,
31'b1100110000000000000010000000000,
31'b0011000000001000000000000100100,
31'b0010000010000000100000100000100,
31'b1100000010000001100000000000000,
31'b0101100000000000000001000001000,
31'b0011000000000000000000000100100,
31'b1001100000000010000000000000001,
31'b1001100000000000000000000000001,
31'b0001000111000000000100000000000,
31'b1100010000000000100000001000000,
31'b0010100000000001001000100000000,
31'b1100100000000000001000000000100,
31'b0000010001000000100010000000000,
31'b1000111000000000000000010000000,
31'b1010100000000000010010000000000,
31'b1000000000000000100001000010000,
31'b0000010100000000000000011000000,
31'b0010000000000000000000101000010,
31'b0010000000000000010000010100000,
31'b0010000000000100000000101000010,
31'b0000010100001000000000011000000,
31'b0011000000100000000000000100100,
31'b1011000000000000000001100000000,
31'b1001100000100000000000000000001,
31'b0000000000001000000000000001100,
31'b0000100100000000010000000010000,
31'b0000000101000001000000010000000,
31'b0001000001000000000000000010100,
31'b0000000000000000000000000001100,
31'b0000000000000010000000000001100,
31'b0000000000000100000000000001100,
31'b0000100000100001000000000000000,
31'b0000000100000000000000101000001,
31'b0000110010001000000000001000000,
31'b0010000001000000100000100000100,
31'b1100000001000001100000000000000,
31'b0000000000010000000000000001100,
31'b0000110010000000000000001000000,
31'b0000000000010100000000000001100,
31'b0000100000110001000000000000000,
31'b0001000100000000000100000000000,
31'b0001000100000010000100000000000,
31'b0001000100000100000100000000000,
31'b0000100000001001000000000000000,
31'b0000000000100000000000000001100,
31'b0000100000000101000000000000000,
31'b0000100000000011000000000000000,
31'b0000100000000001000000000000000,
31'b0001000100010000000100000000000,
31'b1010000000000001000100000000010,
31'b1001000000000010001001000000000,
31'b1001000000000000001001000000000,
31'b0000000000000000001000001000010,
31'b0000100000010101000000000000000,
31'b0000100000010011000000000000000,
31'b0000100000010001000000000000000,
31'b0000000100000101000000010000000,
31'b0001000000000100000000000010100,
31'b0000000100000001000000010000000,
31'b0001000000000000000000000010100,
31'b0000000001000000000000000001100,
31'b0001100000000000000100010000000,
31'b0000000100001001000000010000000,
31'b0001000000001000000000000010100,
31'b0010000000001000000001011000000,
31'b1100000000000101100000000000000,
31'b0010000000000000100000100000100,
31'b1100000000000001100000000000000,
31'b0010000000000000000001011000000,
31'b0011000010000000000000000100100,
31'b0010000000001000100000100000100,
31'b1100000000001001100000000000000,
31'b0001000101000000000100000000000,
31'b0001000101000010000100000000000,
31'b0000100000000000010100000000100,
31'b0001000000100000000000000010100,
31'b0000000000000000010000010010000,
31'b0000100001000101000000000000000,
31'b0000100001000011000000000000000,
31'b0000100001000001000000000000000,
31'b0001010000000000001010000010000,
31'b1100000000000000001010000000010,
31'b0010000010000000010000010100000,
31'b1100000000100001100000000000000,
31'b0000000001000000001000001000010,
31'b0100000000000100001000000010001,
31'b0100000000000010001000000010001,
31'b0100000000000000001000000010001,
31'b1000100000000000000000000000000,
31'b1000100000000010000000000000000,
31'b1000100000000100000000000000000,
31'b1000100000000110000000000000000,
31'b1000100000001000000000000000000,
31'b1000100000001010000000000000000,
31'b1000100000001100000000000000000,
31'b1001000100000001000100000000000,
31'b1000100000010000000000000000000,
31'b1000100000010010000000000000000,
31'b1000100000010100000000000000000,
31'b1000100000010110000000000000000,
31'b0000000000000000000010010100000,
31'b0000001100000000000000001000000,
31'b0010000000000000000100000000010,
31'b0010000000000010000100000000010,
31'b1000100000100000000000000000000,
31'b0100001000000000000000000100000,
31'b1000100000100100000000000000000,
31'b1000000000000001000000000001100,
31'b1000100000101000000000000000000,
31'b1000000101000000000000010000000,
31'b1000100000101100000000000000000,
31'b1000000101000100000000010000000,
31'b1000100000110000000000000000000,
31'b1000000000000000100010001000000,
31'b1000100000110100000000000000000,
31'b1000000000010001000000000001100,
31'b0100000001000000100000000000000,
31'b0100000001000010100000000000000,
31'b0100000001000100100000000000000,
31'b0110001010000000000000000010000,
31'b1000100001000000000000000000000,
31'b1000100001000010000000000000000,
31'b1000100001000100000000000000000,
31'b1000100001000110000000000000000,
31'b1000100001001000000000000000000,
31'b1000000100100000000000010000000,
31'b1000100001001100000000000000000,
31'b1001100000000000000000000011000,
31'b1000100001010000000000000000000,
31'b1100000000000000000000011100000,
31'b1100000000000000010000100000010,
31'b0010010000000000000101000000001,
31'b0100000000100000100000000000000,
31'b0100000000100010100000000000000,
31'b0100000000100100100000000000000,
31'b0100000010000000000000001000110,
31'b1000100001100000000000000000000,
31'b1000000100001000000000010000000,
31'b1000100001100100000000000000000,
31'b1000000100001100000000010000000,
31'b0100000000010000100000000000000,
31'b1000000100000000000000010000000,
31'b1000000000000000010100000001000,
31'b1000000100000100000000010000000,
31'b0100000000001000100000000000000,
31'b0100000000001010100000000000000,
31'b0100000000001100100000000000000,
31'b0101000010000000000000100100000,
31'b0100000000000000100000000000000,
31'b0100000000000010100000000000000,
31'b0100000000000100100000000000000,
31'b0100000000000110100000000000000,
31'b1000100010000000000000000000000,
31'b1000100010000010000000000000000,
31'b1000100010000100000000000000000,
31'b1000100010000110000000000000000,
31'b1000100010001000000000000000000,
31'b1000100010001010000000000000000,
31'b1000100010001100000000000000000,
31'b0100001000000000010001001000000,
31'b1000100010010000000000000000000,
31'b1000100010010010000000000000000,
31'b1000000000000000000010000000110,
31'b1000100000000000101000000001000,
31'b0000000000000000000000000010101,
31'b0000001110000000000000001000000,
31'b0010000010000000000100000000010,
31'b0110001000100000000000000010000,
31'b1000100010100000000000000000000,
31'b1000010000000000001000000000010,
31'b1000100010100100000000000000000,
31'b1000010000000100001000000000010,
31'b1000100010101000000000000000000,
31'b1000010000001000001000000000010,
31'b0101001000000000100000100000000,
31'b0100000001000000001000000001000,
31'b1000100010110000000000000000000,
31'b1000010000010000001000000000010,
31'b1000110000000001000000001000000,
31'b0110001000001000000000000010000,
31'b0100000011000000100000000000000,
31'b0110001000000100000000000010000,
31'b0110001000000010000000000010000,
31'b0110001000000000000000000010000,
31'b1000100011000000000000000000000,
31'b1010010000000000000001010000000,
31'b1000100011000100000000000000000,
31'b0100000000101000001000000001000,
31'b1000100011001000000000000000000,
31'b1010100000000000001000100000000,
31'b0100010000000001100000001000000,
31'b0100000000100000001000000001000,
31'b1101000000000000000001000000100,
31'b0011000000000001000001100000000,
31'b1001101000000000000000100000000,
31'b0001000000000000000000000001101,
31'b0100000010100000100000000000000,
31'b0100000010100010100000000000000,
31'b0100000010100100100000000000000,
31'b0100000000000000000000001000110,
31'b1000100011100000000000000000000,
31'b1000010001000000001000000000010,
31'b0110000000000000100000000110000,
31'b0100000000001000001000000001000,
31'b1000000000000000001001000000001,
31'b1000000110000000000000010000000,
31'b0100000000000010001000000001000,
31'b0100000000000000001000000001000,
31'b0100000010001000100000000000000,
31'b0101000000000100000000100100000,
31'b0101000000000010000000100100000,
31'b0101000000000000000000100100000,
31'b0100000010000000100000000000000,
31'b0100000010000010100000000000000,
31'b0100000010000100100000000000000,
31'b0000000100000000000100000000001,
31'b1000100100000000000000000000000,
31'b1000100100000010000000000000000,
31'b1000100100000100000000000000000,
31'b1001000000001001000100000000000,
31'b1000100100001000000000000000000,
31'b0000001000010000000000001000000,
31'b1001000000000011000100000000000,
31'b1001000000000001000100000000000,
31'b1000100100010000000000000000000,
31'b0000001000001000000000001000000,
31'b1001001000000000000001000000010,
31'b0000100000000000001101000000000,
31'b0000001000000010000000001000000,
31'b0000001000000000000000001000000,
31'b0010000100000000000100000000010,
31'b0000001000000100000000001000000,
31'b1000100100100000000000000000000,
31'b1000000001001000000000010000000,
31'b1001000000000000000000010011000,
31'b1000000100000001000000000001100,
31'b1000000001000010000000010000000,
31'b1000000001000000000000010000000,
31'b1000100000000001010000000010000,
31'b1000000001000100000000010000000,
31'b1000100100110000000000000000000,
31'b0000100001000000000010000100000,
31'b0011000000000000000000000001110,
31'b0000100001000100000010000100000,
31'b0100000101000000100000000000000,
31'b0000001000100000000000001000000,
31'b0110000000000000000000001000101,
31'b0000001000100100000000001000000,
31'b0000000000000000100000001100000,
31'b1000000000101000000000010000000,
31'b1001000000000000010000000000100,
31'b1001000000000010010000000000100,
31'b1000000000100010000000010000000,
31'b1000000000100000000000010000000,
31'b1001000000001000010000000000100,
31'b1000000000100100000000010000000,
31'b1100001000000000000010000000000,
31'b0000100000100000000010000100000,
31'b1100001000000100000010000000000,
31'b0000100001000000001101000000000,
31'b0100000100100000100000000000000,
31'b0000001001000000000000001000000,
31'b0100001000000000000000000010011,
31'b0000001001000100000000001000000,
31'b1000000000001010000000010000000,
31'b1000000000001000000000010000000,
31'b1001000000100000010000000000100,
31'b1000000000001100000000010000000,
31'b1000000000000010000000010000000,
31'b1000000000000000000000010000000,
31'b1000000000000110000000010000000,
31'b1000000000000100000000010000000,
31'b0100000100001000100000000000000,
31'b0000100000000000000010000100000,
31'b0100000100001100100000000000000,
31'b0000100000000100000010000100000,
31'b0100000100000000100000000000000,
31'b1000000000010000000000010000000,
31'b0100000100000100100000000000000,
31'b0000000010000000000100000000001,
31'b1000100110000000000000000000000,
31'b1000100110000010000000000000000,
31'b1101000000000000000010100000000,
31'b0011000000000001000010000000100,
31'b1000100110001000000000000000000,
31'b1000010000000000000000100000001,
31'b0101000000000001011000000000000,
31'b0001000001000000000000101000000,
31'b1000100110010000000000000000000,
31'b0000100000000000010000000001001,
31'b1100100000000000010001000000000,
31'b0000100010000000001101000000000,
31'b0000001010000010000000001000000,
31'b0000001010000000000000001000000,
31'b0010000110000000000100000000010,
31'b0000001010000100000000001000000,
31'b1010000000000000001000110000000,
31'b1000010100000000001000000000010,
31'b0000011000001011000000000000000,
31'b0000011000001001000000000000000,
31'b1010110000000000000001000000000,
31'b1000000011000000000000010000000,
31'b0000011000000011000000000000000,
31'b0000011000000001000000000000000,
31'b0011010000000001001000000000000,
31'b0000100011000000000010000100000,
31'b0000010000000000000101000000010,
31'b0000001000000000010001000100000,
31'b0100000111000000100000000000000,
31'b0000001010100000000000001000000,
31'b0000001000000000100000000000110,
31'b0000000001000000000100000000001,
31'b1000000000000000000001100000010,
31'b1000000010101000000000010000000,
31'b1001000010000000010000000000100,
31'b0001000000001000000000101000000,
31'b1000000010100010000000010000000,
31'b1000000010100000000000010000000,
31'b0001000000000010000000101000000,
31'b0001000000000000000000101000000,
31'b1100001010000000000010000000000,
31'b0000100010100000000010000100000,
31'b0010010000000000001100010000000,
31'b0000000000101000000100000000001,
31'b0110001000000000000100000000100,
31'b0000001011000000000000001000000,
31'b0010000000000000100000001010000,
31'b0000000000100000000100000000001,
31'b1000000010001010000000010000000,
31'b1000000010001000000000010000000,
31'b0000000000001000110001000000000,
31'b0000000000000000000000000100110,
31'b1000000010000010000000010000000,
31'b1000000010000000000000010000000,
31'b0000000000000000110001000000000,
31'b0000000000010000000100000000001,
31'b0101010000000000000110000000000,
31'b0000100010000000000010000100000,
31'b0000010000000001100000000100000,
31'b0000000000001000000100000000001,
31'b0100000110000000100000000000000,
31'b0000000000000100000100000000001,
31'b0000000000000010000100000000001,
31'b0000000000000000000100000000001,
31'b1000101000000000000000000000000,
31'b0100000000100000000000000100000,
31'b1000101000000100000000000000000,
31'b0010000000000001000001000000000,
31'b1000101000001000000000000000000,
31'b0000000100010000000000001000000,
31'b1000101000001100000000000000000,
31'b0010000000001001000001000000000,
31'b1000101000010000000000000000000,
31'b0000000100001000000000001000000,
31'b1001000100000000000001000000010,
31'b0010000000010001000001000000000,
31'b0000000100000010000000001000000,
31'b0000000100000000000000001000000,
31'b0010001000000000000100000000010,
31'b0000000100000100000000001000000,
31'b0100000000000010000000000100000,
31'b0100000000000000000000000100000,
31'b0100000000000110000000000100000,
31'b0100000000000100000000000100000,
31'b0100000000001010000000000100000,
31'b0100000000001000000000000100000,
31'b0101000010000000100000100000000,
31'b0100000000001100000000000100000,
31'b0100000000010010000000000100000,
31'b0100000000010000000000000100000,
31'b0100000001000000001000100010000,
31'b0100000000010100000000000100000,
31'b0100001001000000100000000000000,
31'b0000000100100000000000001000000,
31'b0110000010000010000000000010000,
31'b0110000010000000000000000010000,
31'b1000101001000000000000000000000,
31'b0000000000000000100010010000000,
31'b1000101001000100000000000000000,
31'b0010000001000001000001000000000,
31'b1000101001001000000000000000000,
31'b0000000101010000000000001000000,
31'b0010010000000001000000000000011,
31'b0010000001001001000001000000000,
31'b1100000100000000000010000000000,
31'b0000000101001000000000001000000,
31'b1100000100000100000010000000000,
31'b0010000001010001000001000000000,
31'b0100001000100000100000000000000,
31'b0000000101000000000000001000000,
31'b0100001000100100100000000000000,
31'b0010000000000000100000000000101,
31'b0100000001000010000000000100000,
31'b0100000001000000000000000100000,
31'b0100000001000110000000000100000,
31'b0100000001000100000000000100000,
31'b1000000000000000000010001100000,
31'b1000001100000000000000010000000,
31'b1000001000000000010100000001000,
31'b1000010000000000000000000101010,
31'b0000100000000000000000011000000,
31'b0100000001010000000000000100000,
31'b0100000000000000001000100010000,
31'b0100000001010100000000000100000,
31'b0100001000000000100000000000000,
31'b0100001000000010100000000000000,
31'b0100001000000100100000000000000,
31'b0110000011000000000000000010000,
31'b1000101010000000000000000000000,
31'b0000010000000000010000000010000,
31'b1000101010000100000000000000000,
31'b0010000010000001000001000000000,
31'b1000101010001000000000000000000,
31'b0000010000001000010000000010000,
31'b0101000000100000100000100000000,
31'b0100000000000000010001001000000,
31'b1000101010010000000000000000000,
31'b0000010000010000010000000010000,
31'b1001100001000000000000100000000,
31'b0110000000101000000000000010000,
31'b0000001000000000000000000010101,
31'b0000000110000000000000001000000,
31'b0110000000100010000000000010000,
31'b0110000000100000000000000010000,
31'b0100000010000010000000000100000,
31'b0100000010000000000000000100000,
31'b0101000000001000100000100000000,
31'b0100000010000100000000000100000,
31'b0101000000000100100000100000000,
31'b0100000010001000000000000100000,
31'b0101000000000000100000100000000,
31'b0000010100000001000000000000000,
31'b0111000001000000000000000001000,
31'b0100000010010000000000000100000,
31'b0110000000001010000000000010000,
31'b0110000000001000000000000010000,
31'b0110000000000110000000000010000,
31'b0110000000000100000000000010000,
31'b0110000000000010000000000010000,
31'b0110000000000000000000000010000,
31'b1000101011000000000000000000000,
31'b0000010001000000010000000010000,
31'b1000000000000000010011000000000,
31'b1010100000000000100000000010000,
31'b0011000000000000000100100000010,
31'b0001010100000000000100010000000,
31'b0001010000000000010000000001000,
31'b0100001000100000001000000001000,
31'b1100000110000000000010000000000,
31'b0000010001010000010000000010000,
31'b1001100000000000000000100000000,
31'b1001100000000010000000100000000,
31'b0110000100000000000100000000100,
31'b0000000111000000000000001000000,
31'b1001100000001000000000100000000,
31'b0110000001100000000000000010000,
31'b0111000000010000000000000001000,
31'b0100000011000000000000000100000,
31'b1000100000000000000100001000001,
31'b0100001000001000001000000001000,
31'b1000001000000000001001000000001,
31'b1000001110000000000000010000000,
31'b0101000001000000100000100000000,
31'b0100001000000000001000000001000,
31'b0111000000000000000000000001000,
31'b0111000000000010000000000001000,
31'b1010000000000000000010001010000,
31'b1011000000000000000001000000001,
31'b0100001010000000100000000000000,
31'b0110000001000100000000000010000,
31'b0110000001000010000000000010000,
31'b0110000001000000000000000010000,
31'b1000101100000000000000000000000,
31'b0000000000011000000000001000000,
31'b1001000000010000000001000000010,
31'b0010000100000001000001000000000,
31'b0000000000010010000000001000000,
31'b0000000000010000000000001000000,
31'b0000100000000001001000000000010,
31'b0000000000010100000000001000000,
31'b0000000000001010000000001000000,
31'b0000000000001000000000001000000,
31'b1001000000000000000001000000010,
31'b0000000000001100000000001000000,
31'b0000000000000010000000001000000,
31'b0000000000000000000000001000000,
31'b0000000000000110000000001000000,
31'b0000000000000100000000001000000,
31'b0100000100000010000000000100000,
31'b0100000100000000000000000100000,
31'b0100010000000000000110100000000,
31'b0100000100000100000000000100000,
31'b0000100000000000100010000000000,
31'b0000000000110000000000001000000,
31'b0000100000000100100010000000000,
31'b0000010010000001000000000000000,
31'b1000000000000000100000010100000,
31'b0000000000101000000000001000000,
31'b1001000000100000000001000000010,
31'b0000000010000000010001000100000,
31'b0000000000100010000000001000000,
31'b0000000000100000000000001000000,
31'b0000000010000000100000000000110,
31'b0000000000100100000000001000000,
31'b1100000000010000000010000000000,
31'b0000000100000000100010010000000,
31'b1100000000010100000010000000000,
31'b0010000101000001000001000000000,
31'b0100100000000000000000010100000,
31'b0000000001010000000000001000000,
31'b0100100000000100000000010100000,
31'b0000000001010100000000001000000,
31'b1100000000000000000010000000000,
31'b0000000001001000000000001000000,
31'b1100000000000100000010000000000,
31'b0000000001001100000000001000000,
31'b0000000001000010000000001000000,
31'b0000000001000000000000001000000,
31'b0100000000000000000000000010011,
31'b0000000001000100000000001000000,
31'b1100000000110000000010000000000,
31'b1000001000001000000000010000000,
31'b0011000000000000010001000001000,
31'b1100010000000000001000000000100,
31'b1000001000000010000000010000000,
31'b1000001000000000000000010000000,
31'b1010010000000000010010000000000,
31'b1000001000000100000000010000000,
31'b1100000000100000000010000000000,
31'b0000101000000000000010000100000,
31'b1100000000100100000010000000000,
31'b0000101000000100000010000100000,
31'b0100001100000000100000000000000,
31'b0000000001100000000000001000000,
31'b0100001100000100100000000000000,
31'b0000001010000000000100000000001,
31'b1000101110000000000000000000000,
31'b0000010100000000010000000010000,
31'b0010000000000010000000001110000,
31'b0010000000000000000000001110000,
31'b0000110000000000000000000001100,
31'b0000000010010000000000001000000,
31'b0000010000100011000000000000000,
31'b0000010000100001000000000000000,
31'b1000000000000000010000100000100,
31'b0000000010001000000000001000000,
31'b1001000010000000000001000000010,
31'b0000000010001100000000001000000,
31'b0000000010000010000000001000000,
31'b0000000010000000000000001000000,
31'b0000000010000110000000001000000,
31'b0000000010000100000000001000000,
31'b0101000000000001000010000000001,
31'b0100000110000000000000000100000,
31'b0000010000001011000000000000000,
31'b0000010000001001000000000000000,
31'b0000100010000000100010000000000,
31'b0000010000000101000000000000000,
31'b0000010000000011000000000000000,
31'b0000010000000001000000000000000,
31'b1000000010000000100000010100000,
31'b0000000010101000000000001000000,
31'b0000000000001000100000000000110,
31'b0000000000000000010001000100000,
31'b0000000010100010000000001000000,
31'b0000000010100000000000001000000,
31'b0000000000000000100000000000110,
31'b0000010000010001000000000000000,
31'b1100000010010000000010000000000,
31'b0001010000001000000100010000000,
31'b1100100000000000000000000000110,
31'b0010100000000001000000100000010,
31'b0110000000010000000100000000100,
31'b0001010000000000000100010000000,
31'b0001010100000000010000000001000,
31'b0001001000000000000000101000000,
31'b1100000010000000000010000000000,
31'b0000000011001000000000001000000,
31'b1100000010000100000010000000000,
31'b0000001000101000000100000000001,
31'b0110000000000000000100000000100,
31'b0000000011000000000000001000000,
31'b0110000000000100000100000000100,
31'b0000001000100000000100000000001,
31'b0011000000000000001100000000001,
31'b1100000000000001000000000001010,
31'b0000010000000000010100000000100,
31'b0000010001001001000000000000000,
31'b1000001010000010000000010000000,
31'b1000001010000000000000010000000,
31'b0000010001000011000000000000000,
31'b0000010001000001000000000000000,
31'b1100000010100000000010000000000,
31'b0000101010000000000010000100000,
31'b0000011000000001100000000100000,
31'b0000001000001000000100000000001,
31'b0110000000100000000100000000100,
31'b0000001000000100000100000000001,
31'b0000001000000010000100000000001,
31'b0000001000000000000100000000001,
31'b1000110000000000000000000000000,
31'b1000110000000010000000000000000,
31'b1000110000000100000000000000000,
31'b1000110000000110000000000000000,
31'b1000110000001000000000000000000,
31'b1000110000001010000000000000000,
31'b1100000000000000100100100000000,
31'b0010001000010000010000000100000,
31'b1000110000010000000000000000000,
31'b1000110000010010000000000000000,
31'b1000110000010100000000000000000,
31'b0101000000000000000000010100001,
31'b0000000000000000010000100001000,
31'b0000011100000000000000001000000,
31'b0010010000000000000100000000010,
31'b0010001000000000010000000100000,
31'b1000110000100000000000000000000,
31'b1000000010000000001000000000010,
31'b1000110000100100000000000000000,
31'b1000010000000001000000000001100,
31'b1010000001000000000000100000010,
31'b1000010101000000000000010000000,
31'b0001001000000000000010000100001,
31'b0000001110000001000000000000000,
31'b1000110000110000000000000000000,
31'b1000010000000000100010001000000,
31'b1000000000000000100000000001010,
31'b1000100000000000001010000000100,
31'b0100010001000000100000000000000,
31'b0100010001000010100000000000000,
31'b1110100000000000010000000000000,
31'b0010100010000000001100000000000,
31'b1000110001000000000000000000000,
31'b1010000010000000000001010000000,
31'b0010000000000000110000000000000,
31'b0010000000000010110000000000000,
31'b1010000000100000000000100000010,
31'b1000100000000000000001000000011,
31'b0100100000000000000000000001010,
31'b0100100000000010000000000001010,
31'b1110000000000000000100000001000,
31'b0010000010000000011000000001000,
31'b0010000000010000110000000000000,
31'b0010000000000000000101000000001,
31'b0100010000100000100000000000000,
31'b0100010000100010100000000000000,
31'b0100100000010000000000000001010,
31'b1001001100000000000000000000001,
31'b1010000000001000000000100000010,
31'b1000010100001000000000010000000,
31'b0010000000100000110000000000000,
31'b0011000000000000000001101000000,
31'b1010000000000000000000100000010,
31'b1000010100000000000000010000000,
31'b1010000000000100000000100000010,
31'b1000010100000100000000010000000,
31'b0100010000001000100000000000000,
31'b0100010000001010100000000000000,
31'b0000100000000000000100100000000,
31'b0001000000000000100010000000001,
31'b0100010000000000100000000000000,
31'b0100010000000010100000000000000,
31'b0100010000000100100000000000000,
31'b0100100010000001000010000000000,
31'b1000110010000000000000000000000,
31'b0000001000000000010000000010000,
31'b1000110010000100000000000000000,
31'b1000000000000001100010000000000,
31'b1000110010001000000000000000000,
31'b1000000100000000000000100000001,
31'b0100000100000000000001100001000,
31'b0000001100100001000000000000000,
31'b1000110010010000000000000000000,
31'b1000000000000000000000001001100,
31'b1000100000100001000000001000000,
31'b1000000000010001100010000000000,
31'b0000010000000000000000000010101,
31'b1000000100010000000000100000001,
31'b0011000000000000011000000010000,
31'b0010100000100000001100000000000,
31'b1000000000000010001000000000010,
31'b1000000000000000001000000000010,
31'b1000100000010001000000001000000,
31'b1000000000000100001000000000010,
31'b1010100100000000000001000000000,
31'b1000000000001000001000000000010,
31'b0001000000000000001001001000000,
31'b0000001100000001000000000000000,
31'b1000100000000101000000001000000,
31'b1000000000010000001000000000010,
31'b1000100000000001000000001000000,
31'b1000100000000011000000001000000,
31'b0100010011000000100000000000000,
31'b1001000100000000000100001000000,
31'b1011001000000000000000000000010,
31'b0010100000000000001100000000000,
31'b1010000000000010000001010000000,
31'b1010000000000000000001010000000,
31'b0010000010000000110000000000000,
31'b1010000000000100000001010000000,
31'b0100000000010000000010000001100,
31'b1010000000001000000001010000000,
31'b0100000000000001100000001000000,
31'b0100010000100000001000000001000,
31'b0110000100000000100001000000000,
31'b0010000000000000011000000001000,
31'b0010000100000000001100010000000,
31'b0010000010000000000101000000001,
31'b0100000000000000000010000001100,
31'b0100100000000000101000000000010,
31'b1001000000000000000000001010100,
31'b1000000100000001000000011000000,
31'b1000100000000000000000110000001,
31'b1000000001000000001000000000010,
31'b0010000010100000110000000000000,
31'b1100000000000001000000010100000,
31'b1010000010000000000000100000010,
31'b1000010110000000000000010000000,
31'b0100010000000010001000000001000,
31'b0100010000000000001000000001000,
31'b0101000100000000000110000000000,
31'b1000000001010000001000000000010,
31'b0000100010000000000100100000000,
31'b0101010000000000000000100100000,
31'b0100010010000000100000000000000,
31'b0100100000000101000010000000000,
31'b0100100000000011000010000000000,
31'b0100100000000001000010000000000,
31'b1000110100000000000000000000000,
31'b1000110100000010000000000000000,
31'b1001000000000000100000000100001,
31'b0100001000010000000001000010000,
31'b1000110100001000000000000000000,
31'b1000000010000000000000100000001,
31'b0100000010000000000001100001000,
31'b0000001010100001000000000000000,
31'b1000110100010000000000000000000,
31'b0000100000000000000000100010100,
31'b0100001000000010000001000010000,
31'b0100001000000000000001000010000,
31'b0000011000000010000000001000000,
31'b0000011000000000000000001000000,
31'b0000001000000000000010000001010,
31'b0000000000000000000100110000000,
31'b1000110100100000000000000000000,
31'b1000010001001000000000010000000,
31'b0100001000000000000110100000000,
31'b0100000000000000000000010001010,
31'b1010100010000000000001000000000,
31'b1000010001000000000000010000000,
31'b0000001010000011000000000000000,
31'b0000001010000001000000000000000,
31'b0011000010000001001000000000000,
31'b0011000000000000000010001000100,
31'b0000000010000000000101000000010,
31'b0100001000100000000001000010000,
31'b0101000000000000011000001000000,
31'b0001000001000001000000100000000,
31'b0000001010010011000000000000000,
31'b0000001010010001000000000000000,
31'b1010000000000000001000000000001,
31'b1010000000000010001000000000001,
31'b0010000100000000110000000000000,
31'b0110000000000000001001000001000,
31'b1010000000001000001000000000001,
31'b1000010000100000000000010000000,
31'b0100100100000000000000000001010,
31'b1001001000010000000000000000001,
31'b1100011000000000000010000000000,
31'b0001001000000000000010000010010,
31'b0010000100010000110000000000000,
31'b1110000000000000010000010000000,
31'b0101001000000000000001000001000,
31'b0001000000100001000000100000000,
31'b1001001000000010000000000000001,
31'b1001001000000000000000000000001,
31'b1010000000100000001000000000001,
31'b1000010000001000000000010000000,
31'b0010001000000001001000100000000,
31'b1100001000000000001000000000100,
31'b1000010000000010000000010000000,
31'b1000010000000000000000010000000,
31'b1010001000000000010010000000000,
31'b1000010000000100000000010000000,
31'b0101000010000000000110000000000,
31'b0001000000001001000000100000000,
31'b0000100100000000000100100000000,
31'b0001000100000000100010000000001,
31'b0100010100000000100000000000000,
31'b0001000000000001000000100000000,
31'b0101100000000000000000000100001,
31'b0001000000000101000000100000000,
31'b1000110110000000000000000000000,
31'b1000000000001000000000100000001,
31'b0100000000010001000010010000000,
31'b0000001000101001000000000000000,
31'b1000000000000010000000100000001,
31'b1000000000000000000000100000001,
31'b0100000000000000000001100001000,
31'b0000001000100001000000000000000,
31'b0110000001000000100001000000000,
31'b1000000100000000000000001001100,
31'b0100000000000001000010010000000,
31'b0100001010000000000001000010000,
31'b1000100000000000010000001010000,
31'b1000000000010000000000100000001,
31'b0100000000010000000001100001000,
31'b0000001000110001000000000000000,
31'b1010100000001000000001000000000,
31'b1000000100000000001000000000010,
31'b0000001000001011000000000000000,
31'b0000001000001001000000000000000,
31'b1010100000000000000001000000000,
31'b0000001000000101000000000000000,
31'b0000001000000011000000000000000,
31'b0000001000000001000000000000000,
31'b0011000000000001001000000000000,
31'b1001000000001000000100001000000,
31'b0000000000000000000101000000010,
31'b0000001000011001000000000000000,
31'b1010100000010000000001000000000,
31'b1001000000000000000100001000000,
31'b0000001000010011000000000000000,
31'b0000001000010001000000000000000,
31'b1010000010000000001000000000001,
31'b1010000100000000000001010000000,
31'b0010000110000000110000000000000,
31'b0001101000000000000000000010100,
31'b1000100000000000001000010000010,
31'b1000000001000000000000100000001,
31'b0100000100000001100000001000000,
31'b0001010000000000000000101000000,
31'b0110000000000000100001000000000,
31'b0110000000000010100001000000000,
31'b0010000000000000001100010000000,
31'b1010000000000000100000000001001,
31'b0110000000001000100001000000000,
31'b1000000001010000000000100000001,
31'b1000000000000011000000011000000,
31'b1000000000000001000000011000000,
31'b0101000000010000000110000000000,
31'b1000010010001000000000010000000,
31'b0000001000000000010100000000100,
31'b0000010000000000000000000100110,
31'b1010100001000000000001000000000,
31'b1000010010000000000000010000000,
31'b0000010000000000110001000000000,
31'b0000001001000001000000000000000,
31'b0101000000000000000110000000000,
31'b0101000000000010000110000000000,
31'b0000000000000001100000000100000,
31'b0000010000001000000100000000001,
31'b0101000000001000000110000000000,
31'b0001000010000001000000100000000,
31'b0000010000000010000100000000001,
31'b0000010000000000000100000000001,
31'b1000111000000000000000000000000,
31'b0000000010000000010000000010000,
31'b1000111000000100000000000000000,
31'b0010010000000001000001000000000,
31'b1000111000001000000000000000000,
31'b0000010100010000000000001000000,
31'b0010000001000001000000000000011,
31'b0010000000010000010000000100000,
31'b1000111000010000000000000000000,
31'b0000010100001000000000001000000,
31'b0100000100000010000001000010000,
31'b0100000100000000000001000010000,
31'b0000010100000010000000001000000,
31'b0000010100000000000000001000000,
31'b0010000000000010010000000100000,
31'b0010000000000000010000000100000,
31'b0100010000000010000000000100000,
31'b0100010000000000000000000100000,
31'b0100010000000110000000000100000,
31'b0100010000000100000000000100000,
31'b0100010000001010000000000100000,
31'b0100010000001000000000000100000,
31'b0001000000000000000010000100001,
31'b0000000110000001000000000000000,
31'b0100010000010010000000000100000,
31'b0100010000010000000000000100000,
31'b1001100000000000000000010000001,
31'b0100010000010100000000000100000,
31'b0100011001000000100000000000000,
31'b0100000000000001010001000000000,
31'b1011000010000000000000000000010,
31'b0010000000100000010000000100000,
31'b1010000000000001000010000010000,
31'b0000010000000000100010010000000,
31'b0010001000000000110000000000000,
31'b0010010001000001000001000000000,
31'b0010000000000101000000000000011,
31'b0001000110000000000100010000000,
31'b0010000000000001000000000000011,
31'b1001000100010000000000000000001,
31'b1100010100000000000010000000000,
31'b0001000100000000000010000010010,
31'b0010001000010000110000000000000,
31'b1100000000000000000100100100000,
31'b0101000100000000000001000001000,
31'b0001000000000000111000000000000,
31'b1001000100000010000000000000001,
31'b1001000100000000000000000000001,
31'b0100010001000010000000000100000,
31'b0100010001000000000000000100000,
31'b0010001000100000110000000000000,
31'b1100000100000000001000000000100,
31'b1010001000000000000000100000010,
31'b1000011100000000000000010000000,
31'b1010000100000000010010000000000,
31'b1000000000000000000000000101010,
31'b0100000000000000000101000000100,
31'b0100010001010000000000000100000,
31'b0000101000000000000100100000000,
31'b1001000000000000001000100000010,
31'b0100011000000000100000000000000,
31'b0100011000000010100000000000000,
31'b0100100000000000000001010010000,
31'b1001000100100000000000000000001,
31'b0000000000000010010000000010000,
31'b0000000000000000010000000010000,
31'b0000100001000001000000010000000,
31'b0000000000000100010000000010000,
31'b0000100100000000000000000001100,
31'b0000000000001000010000000010000,
31'b0001000001000000010000000001000,
31'b0000000100100001000000000000000,
31'b0000100000000000000000101000001,
31'b0000000000010000010000000010000,
31'b0100000000000011000000001100000,
31'b0100000000000001000000001100000,
31'b0000100100010000000000000001100,
31'b0000010110000000000000001000000,
31'b1011000000100000000000000000010,
31'b0010000010000000010000000100000,
31'b0001100000000000000100000000000,
31'b0000000000100000010000000010000,
31'b0001100000000100000100000000000,
31'b0000000100001001000000000000000,
31'b0001100000001000000100000000000,
31'b0000000100000101000000000000000,
31'b0000000100000011000000000000000,
31'b0000000100000001000000000000000,
31'b0010000000000010000001001000000,
31'b0010000000000000000001001000000,
31'b1011000000001000000000000000010,
31'b0010000000000100000001001000000,
31'b1011000000000100000000000000010,
31'b0010000000001000000001001000000,
31'b1011000000000000000000000000010,
31'b0000000100010001000000000000000,
31'b0000100000000101000000010000000,
31'b0000000001000000010000000010000,
31'b0000100000000001000000010000000,
31'b0000100000000011000000010000000,
31'b0001000000000100010000000001000,
31'b0001000100000000000100010000000,
31'b0001000000000000010000000001000,
31'b0001000000000010010000000001000,
31'b0000100001000000000000101000001,
31'b0000000001010000010000000010000,
31'b0000100000010001000000010000000,
31'b0100100000000000000000100010010,
31'b1101000000000000100100000000000,
31'b0001000100010000000100010000000,
31'b1000000000000001000010000100000,
31'b1001000110000000000000000000001,
31'b0001100001000000000100000000000,
31'b0000000000000000000000010001100,
31'b0000100000100001000000010000000,
31'b0000000101001001000000000000000,
31'b0001100001001000000100000000000,
31'b0000000101000101000000000000000,
31'b0001000000100000010000000001000,
31'b0000000101000001000000000000000,
31'b0111010000000000000000000001000,
31'b0010000001000000000001001000000,
31'b0000101010000000000100100000000,
31'b0010000001000100000001001000000,
31'b1110000000000000000011000000000,
31'b0010000001001000000001001000000,
31'b1011000001000000000000000000010,
31'b0010000000000000000010000001001,
31'b1000111100000000000000000000000,
31'b0000010000011000000000001000000,
31'b0100000000100000000110100000000,
31'b0100000000010000000001000010000,
31'b0000100010000000000000000001100,
31'b0000010000010000000000001000000,
31'b0000000010100011000000000000000,
31'b0000000010100001000000000000000,
31'b1000000000000000000000000011001,
31'b0000010000001000000000001000000,
31'b0100000000000010000001000010000,
31'b0100000000000000000001000010000,
31'b0000010000000010000000001000000,
31'b0000010000000000000000001000000,
31'b0000000000000000000010000001010,
31'b0000010000000100000000001000000,
31'b0100010100000010000000000100000,
31'b0100010100000000000000000100000,
31'b0100000000000000000110100000000,
31'b0000000010001001000000000000000,
31'b0000110000000000100010000000000,
31'b0000000010000101000000000000000,
31'b0000000010000011000000000000000,
31'b0000000010000001000000000000000,
31'b1000010000000000100000010100000,
31'b0010000000000001000000000110000,
31'b0100000000100010000001000010000,
31'b0100000000100000000001000010000,
31'b0000010000100010000000001000000,
31'b0000010000100000000000001000000,
31'b0000000010010011000000000000000,
31'b0000000010010001000000000000000,
31'b1100010000010000000010000000000,
31'b0001000010001000000100010000000,
31'b0010001100000000110000000000000,
31'b1100000000100000001000000000100,
31'b0101000000010000000001000001000,
31'b0001000010000000000100010000000,
31'b1010000000100000010010000000000,
31'b1001000000010000000000000000001,
31'b1100010000000000000010000000000,
31'b0001000000000000000010000010010,
31'b1100010000000100000010000000000,
31'b1001000000001000000000000000001,
31'b0101000000000000000001000001000,
31'b0000010001000000000000001000000,
31'b1001000000000010000000000000001,
31'b1001000000000000000000000000001,
31'b0010000000000101001000100000000,
31'b1100000000000100001000000000100,
31'b0010000000000001001000100000000,
31'b1100000000000000001000000000100,
31'b1010000000000100010010000000000,
31'b1000011000000000000000010000000,
31'b1010000000000000010010000000000,
31'b0000000011000001000000000000000,
31'b1100010000100000000010000000000,
31'b0010100000000000000000101000010,
31'b0010100000000000010000010100000,
31'b1100000000010000001000000000100,
31'b0101000000100000000001000001000,
31'b0001001000000001000000100000000,
31'b1010000000010000010010000000000,
31'b1001000000100000000000000000001,
31'b0000100000001000000000000001100,
31'b0000000100000000010000000010000,
31'b0000000000101011000000000000000,
31'b0000000000101001000000000000000,
31'b0000100000000000000000000001100,
31'b0000000000100101000000000000000,
31'b0000000000100011000000000000000,
31'b0000000000100001000000000000000,
31'b1000010000000000010000100000100,
31'b0000010010001000000000001000000,
31'b0100001000000001000010010000000,
31'b0100000010000000000001000010000,
31'b0000100000010000000000000001100,
31'b0000010010000000000000001000000,
31'b0000000010000000000010000001010,
31'b0000000000110001000000000000000,
31'b0001100100000000000100000000000,
31'b0000000000001101000000000000000,
31'b0000000000001011000000000000000,
31'b0000000000001001000000000000000,
31'b0000000000000111000000000000000,
31'b0000000000000101000000000000000,
31'b0000000000000011000000000000000,
31'b0000000000000001000000000000000,
31'b0011001000000001001000000000000,
31'b0010000100000000000001001000000,
31'b0000001000000000000101000000010,
31'b0000000000011001000000000000000,
31'b0000100000000000001000001000010,
31'b0000000000010101000000000000000,
31'b0000000000010011000000000000000,
31'b0000000000010001000000000000000,
31'b0001000000100001000000000011000,
31'b0001000000001000000100010000000,
31'b0000100100000001000000010000000,
31'b0001100000000000000000000010100,
31'b0001000000000010000100010000000,
31'b0001000000000000000100010000000,
31'b0001000100000000010000000001000,
31'b0000000001100001000000000000000,
31'b1100010010000000000010000000000,
31'b0001000010000000000010000010010,
31'b0010100000000000100000100000100,
31'b1100100000000001100000000000000,
31'b0110010000000000000100000000100,
31'b0001000000010000000100010000000,
31'b1001000010000010000000000000001,
31'b1001000010000000000000000000001,
31'b0001000000000001000000000011000,
31'b0000000100000000000000010001100,
31'b0000000000000000010100000000100,
31'b0000000001001001000000000000000,
31'b0000100000000000010000010010000,
31'b0000000001000101000000000000000,
31'b0000000001000011000000000000000,
31'b0000000001000001000000000000000,
31'b1100000000000000100000000001100,
31'b0010000101000000000001001000000,
31'b0000001000000001100000000100000,
31'b0000000001011001000000000000000,
31'b0000100001000000001000001000010,
31'b0000000001010101000000000000000,
31'b0000000001010011000000000000000,
31'b0000000001010001000000000000000,
31'b1001000000000000000000000000000,
31'b1001000000000010000000000000000,
31'b1001000000000100000000000000000,
31'b1001000000000110000000000000000,
31'b1001000000001000000000000000000,
31'b1001000000001010000000000000000,
31'b1001000000001100000000000000000,
31'b0000000000000000000001001000010,
31'b1001000000010000000000000000000,
31'b1001000000010010000000000000000,
31'b1001000000010100000000000000000,
31'b1010001000001000001000000000000,
31'b1001000000011000000000000000000,
31'b1010001000000100001000000000000,
31'b1010001000000010001000000000000,
31'b1010001000000000001000000000000,
31'b1001000000100000000000000000000,
31'b1001000000100010000000000000000,
31'b1001000000100100000000000000000,
31'b1001000000100110000000000000000,
31'b1001000000101000000000000000000,
31'b1001000000101010000000000000000,
31'b1001000000101100000000000000000,
31'b1000000000000000010000010000100,
31'b1001000000110000000000000000000,
31'b1010000000000000010010000000001,
31'b1001000000110100000000000000000,
31'b0100100000000000100000000011000,
31'b1100000000000000001000000000101,
31'b0010000000000100010000000010010,
31'b0110100000000000001000000100000,
31'b0010000000000000010000000010010,
31'b1001000001000000000000000000000,
31'b1001000001000010000000000000000,
31'b0000010000000000000000001000001,
31'b1000000000001000000000000011000,
31'b1001000001001000000000000000000,
31'b1000000000000100000000000011000,
31'b1000000000000010000000000011000,
31'b1000000000000000000000000011000,
31'b1001000001010000000000000000000,
31'b1010000010000000000000000101000,
31'b1000001010000000000000100000000,
31'b1000001010000010000000100000000,
31'b1001000001011000000000000000000,
31'b1001001000000000100000000100000,
31'b1000001010001000000000100000000,
31'b1000000000010000000000000011000,
31'b1001000001100000000000000000000,
31'b1001000001100010000000000000000,
31'b1000000000000001000100010000000,
31'b1000000000101000000000000011000,
31'b1001000001101000000000000000000,
31'b1001100100000000000000010000000,
31'b1000000000100010000000000011000,
31'b1000000000100000000000000011000,
31'b0000000010000001000000000000001,
31'b0001000100000000000010000100000,
31'b0001010000000000000100100000000,
31'b0100100010000000000000100100000,
31'b0101100000000000100000000000000,
31'b0101100000000010100000000000000,
31'b0101100000000100100000000000000,
31'b1000001000000000000001010000010,
31'b1001000010000000000000000000000,
31'b1001000010000010000000000000000,
31'b1001000010000100000000000000000,
31'b1001000010000110000000000000000,
31'b1001000010001000000000000000000,
31'b1001000010001010000000000000000,
31'b1001000010001100000000000000000,
31'b1000000000000000100000100100000,
31'b1001000010010000000000000000000,
31'b1010000001000000000000000101000,
31'b1000001001000000000000100000000,
31'b1001000000000000101000000001000,
31'b1001000010011000000000000000000,
31'b0100010000000000000110010000000,
31'b1011000000000000000000000110000,
31'b1010001010000000001000000000000,
31'b0000011000000000000100000000000,
31'b0000000000000000010000000100010,
31'b0000000000000000000000111000000,
31'b0000000000000100010000000100010,
31'b0000000000000000100001000000100,
31'b0000000000001000010000000100010,
31'b0000000000001000000000111000000,
31'b1000000010000000010000010000100,
31'b0000000001000001000000000000001,
31'b0000000001000011000000000000001,
31'b0000000001000101000000000000001,
31'b0100100001000000000000100100000,
31'b0000000001001001000000000000001,
31'b0000010000000001000001000000010,
31'b0000000101000000100010100000000,
31'b0011010000000000001100000000000,
31'b1001000011000000000000000000000,
31'b1010000000010000000000000101000,
31'b1000001000010000000000100000000,
31'b1000001000010010000000100000000,
31'b1001000011001000000000000000000,
31'b1011000000000000001000100000000,
31'b1000001000011000000000100000000,
31'b1000000010000000000000000011000,
31'b0000000000100001000000000000001,
31'b1010000000000000000000000101000,
31'b1000001000000000000000100000000,
31'b1000001000000010000000100000000,
31'b1000000000000000101000000010000,
31'b1010000000001000000000000101000,
31'b1000001000001000000000100000000,
31'b1000001000001010000000100000000,
31'b0000000000010001000000000000001,
31'b0000000001000000010000000100010,
31'b0000000001000000000000111000000,
31'b0100100000010000000000100100000,
31'b0000000001000000100001000000100,
31'b0000011000000001010000000000100,
31'b0010000100000000000001001000001,
31'b1100000000000000000010110000000,
31'b0000000000000001000000000000001,
31'b0000000000000011000000000000001,
31'b0000000000000101000000000000001,
31'b0100100000000000000000100100000,
31'b0000000000001001000000000000001,
31'b0000010000000000100100000100000,
31'b0000000100000000100010100000000,
31'b0101010000000001000010000000000,
31'b1001000100000000000000000000000,
31'b1001000100000010000000000000000,
31'b1001000100000100000000000000000,
31'b1001000100000110000000000000000,
31'b1001000100001000000000000000000,
31'b1001000100001010000000000000000,
31'b1001000100001100000000000000000,
31'b1000100000000001000100000000000,
31'b1001000100010000000000000000000,
31'b0010000000000001000000000000010,
31'b1001000100010100000000000000000,
31'b0010000000000101000000000000010,
31'b1001000100011000000000000000000,
31'b0010000000001001000000000000010,
31'b0100000010000000000000110100000,
31'b1010001100000000001000000000000,
31'b1001000100100000000000000000000,
31'b1001000100100010000000000000000,
31'b1001000100100100000000000000000,
31'b0100011000000000100000000000001,
31'b1000000000000000000100000001100,
31'b1001100001000000000000010000000,
31'b1001000000000001010000000010000,
31'b1000100000100001000100000000000,
31'b1001000100110000000000000000000,
31'b0010000000100001000000000000010,
31'b0100000000001000110000000000100,
31'b0100000000000000000001000100010,
31'b1101000000000000000000001100000,
31'b0010001000000000000010100010000,
31'b0100000000000000110000000000100,
31'b0100000000001000000001000100010,
31'b1001000101000000000000000000000,
31'b1001000101000010000000000000000,
31'b1000100000000000010000000000100,
31'b1000100000000010010000000000100,
31'b1001000101001000000000000000000,
31'b1001100000100000000000010000000,
31'b1000100000001000010000000000100,
31'b1000000100000000000000000011000,
31'b1001000101010000000000000000000,
31'b0010000001000001000000000000010,
31'b1000100000010000010000000000100,
31'b0110000000000000001000010100000,
31'b0010010000000001000001000000001,
31'b0010011000000000000000000100100,
31'b0000010000000000000000100001100,
31'b1000111000000000000000000000001,
31'b1001000101100000000000000000000,
31'b1000000000000001010000000001000,
31'b1000100000100000010000000000100,
31'b1001000000000000000100000010100,
31'b1001100000000010000000010000000,
31'b1001100000000000000000010000000,
31'b0100010000010000000000000100001,
31'b1001100000000100000000010000000,
31'b0001000000000010000010000100000,
31'b0001000000000000000010000100000,
31'b0100010000001000000000000100001,
31'b0100000000000001100100000000000,
31'b0101100100000000100000000000000,
31'b0001000000001000000010000100000,
31'b0100010000000000000000000100001,
31'b0100010000000010000000000100001,
31'b1001000110000000000000000000000,
31'b1001000110000010000000000000000,
31'b1100100000000000000010100000000,
31'b0010100000000001000010000000100,
31'b1001000110001000000000000000000,
31'b0100000001000000001000010010000,
31'b0100100000000001011000000000000,
31'b0000100001000000000000101000000,
31'b1001000110010000000000000000000,
31'b0010000010000001000000000000010,
31'b1101000000000000010001000000000,
31'b0010010000000000001000000001100,
31'b0100000000000100000000110100000,
31'b0100000000000000010000001000010,
31'b0100000000000000000000110100000,
31'b0100000000000100010000001000010,
31'b0010000000000000000010000001000,
31'b0010000000000010000010000001000,
31'b0010000000000100000010000001000,
31'b0010010000000000000000001000010,
31'b0010000000001000000010000001000,
31'b0110000000000000000001000010010,
31'b0010000001000000000001001000001,
31'b0011000001000000000010000010000,
31'b0010000000010000000010000001000,
31'b0010000010100001000000000000010,
31'b0010000000010100000010000001000,
31'b1100000000000000100000101000000,
31'b0010000000011000000010000001000,
31'b1100000000000000000001010000100,
31'b0000000001000000100010100000000,
31'b1000101000000000000000110000000,
31'b1001000111000000000000000000000,
31'b0100010000000000100100001000000,
31'b1000100010000000010000000000100,
31'b0000100000001000000000101000000,
31'b0100000000000010001000010010000,
31'b0100000000000000001000010010000,
31'b0000100000000010000000101000000,
31'b0000100000000000000000101000000,
31'b1000000000000000010010000000010,
31'b1010000100000000000000000101000,
31'b1000001100000000000000100000000,
31'b1000010000000000010000001001000,
31'b0000000000000100010000000010001,
31'b0100000001000000010000001000010,
31'b0000000000000000010000000010001,
31'b0000100000010000000000101000000,
31'b0010000001000000000010000001000,
31'b1011000000000000000000000000011,
31'b0010000001000100000010000001000,
31'b0011000000001000000010000010000,
31'b0010000001001000000010000001000,
31'b1110000000000000000000001001000,
31'b0010000000000000000001001000001,
31'b0011000000000000000010000010000,
31'b0000000100000001000000000000001,
31'b0001000010000000000010000100000,
31'b0000000100000101000000000000001,
31'b0100100100000000000000100100000,
31'b0000000100001001000000000000001,
31'b0001100000000100000100000000001,
31'b0000000000000000100010100000000,
31'b0001100000000000000100000000001,
31'b1001001000000000000000000000000,
31'b1001001000000010000000000000000,
31'b1001001000000100000000000000000,
31'b1010000000011000001000000000000,
31'b1001001000001000000000000000000,
31'b1010000000010100001000000000000,
31'b1010000000010010001000000000000,
31'b1010000000010000001000000000000,
31'b1001001000010000000000000000000,
31'b1010000000001100001000000000000,
31'b0000000000000001000100001000000,
31'b1010000000001000001000000000000,
31'b1010000000000110001000000000000,
31'b1010000000000100001000000000000,
31'b1010000000000010001000000000000,
31'b1010000000000000001000000000000,
31'b0000010010000000000100000000000,
31'b0101100000000000000000000100000,
31'b0001000000000001000000100000001,
31'b0101100000000100000000000100000,
31'b0001000100000000100010000000000,
31'b0101100000001000000000000100000,
31'b0100100010000000100000100000000,
31'b1010000000110000001000000000000,
31'b0001000001000000000000011000000,
31'b0101100000010000000000000100000,
31'b1000010000000000000000010000001,
31'b1010000000101000001000000000000,
31'b0001000100010000100010000000000,
31'b1101000000000000000010010000000,
31'b1010000000100010001000000000000,
31'b1010000000100000001000000000000,
31'b1001001001000000000000000000000,
31'b1001001001000010000000000000000,
31'b1000000010010000000000100000000,
31'b1000001000001000000000000011000,
31'b1010000000000000000000100110000,
31'b1001000000010000100000000100000,
31'b1000001000000010000000000011000,
31'b1000001000000000000000000011000,
31'b1000000010000100000000100000000,
31'b1001000000001000100000000100000,
31'b1000000010000000000000100000000,
31'b1000000010000010000000100000000,
31'b1001000000000010100000000100000,
31'b1001000000000000100000000100000,
31'b1000000010001000000000100000000,
31'b0000000000000000010000001000100,
31'b0001000000010000000000011000000,
31'b0110010000000000000000001000100,
31'b1000001000000001000100010000000,
31'b0110100000000000101000000000000,
31'b0001000101000000100010000000000,
31'b0010010000000000001100100000000,
31'b0100100000000000000000000111000,
31'b0010000000000000000001000010100,
31'b0001000000000000000000011000000,
31'b0001000000000010000000011000000,
31'b1000000010100000000000100000000,
31'b1000000010100010000000100000000,
31'b0001000000001000000000011000000,
31'b1001000000100000100000000100000,
31'b1000000010101000000000100000000,
31'b1000000000000000000001010000010,
31'b0000010000100000000100000000000,
31'b1000000000000000001000000110000,
31'b1000000001010000000000100000000,
31'b1000000001010010000000100000000,
31'b1010000000000000100000000001000,
31'b1010000000000010100000000001000,
31'b1010000000000100100000000001000,
31'b1010000010010000001000000000000,
31'b1000000001000100000000100000000,
31'b1000000001000110000000100000000,
31'b1000000001000000000000100000000,
31'b1000000001000010000000100000000,
31'b1010000000010000100000000001000,
31'b1010000010000100001000000000000,
31'b1000000001001000000000100000000,
31'b1010000010000000001000000000000,
31'b0000010000000000000100000000000,
31'b0000010000000010000100000000000,
31'b0000010000000100000100000000000,
31'b0000010000000110000100000000000,
31'b0000010000001000000100000000000,
31'b0000010000001010000100000000000,
31'b0100100000000000100000100000000,
31'b0101000000000000000110000000001,
31'b0000010000010000000100000000000,
31'b0000010000010010000100000000000,
31'b1000000001100000000000100000000,
31'b1000010100000000001001000000000,
31'b0000010000011000000100000000000,
31'b0000011000000001000001000000010,
31'b1010110000000000000000000000010,
31'b1010000010100000001000000000000,
31'b1000000000010100000000100000000,
31'b1000000001000000001000000110000,
31'b1000000000010000000000100000000,
31'b1000000000010010000000100000000,
31'b1010000001000000100000000001000,
31'b0100000100000000000001001000100,
31'b1000000000011000000000100000000,
31'b1000001010000000000000000011000,
31'b1000000000000100000000100000000,
31'b1000000000000110000000100000000,
31'b1000000000000000000000100000000,
31'b1000000000000010000000100000000,
31'b1000000000001100000000100000000,
31'b1001000010000000100000000100000,
31'b1000000000001000000000100000000,
31'b1000000000001010000000100000000,
31'b0000010001000000000100000000000,
31'b0000010001000010000100000000000,
31'b1000000000110000000000100000000,
31'b1000000000110010000000100000000,
31'b0000010001001000000100000000000,
31'b0000010000000001010000000000100,
31'b1100000000000000000100000001010,
31'b0011000000000001001000000000001,
31'b0000001000000001000000000000001,
31'b0000000000000000000001000100100,
31'b1000000000100000000000100000000,
31'b1000000000100010000000100000000,
31'b0000000000000000110000000000010,
31'b0000000000001000000001000100100,
31'b1000000000101000000000100000000,
31'b1000000010000000000001010000010,
31'b1001001100000000000000000000000,
31'b1001001100000010000000000000000,
31'b1001001100000100000000000000000,
31'b0100010000100000100000000000001,
31'b0010000000000000000101000000000,
31'b0010000000000010000101000000000,
31'b0010000000000100000101000000000,
31'b1010000100010000001000000000000,
31'b1001001100010000000000000000000,
31'b0010001000000001000000000000010,
31'b1000100000000000000001000000010,
31'b1010000100001000001000000000000,
31'b0010000000010000000101000000000,
31'b0001100000000000000000001000000,
31'b1010000100000010001000000000000,
31'b1010000100000000001000000000000,
31'b0001000000001000100010000000000,
31'b0101100100000000000000000100000,
31'b0100010000000010100000000000001,
31'b0100010000000000100000000000001,
31'b0001000000000000100010000000000,
31'b0001000000000010100010000000000,
31'b0100000000000001000100000100000,
31'b0100010000001000100000000000001,
31'b0001000101000000000000011000000,
31'b0010001000100001000000000000010,
31'b1000100000100000000001000000010,
31'b1010000000000000000000100000011,
31'b0001000000010000100010000000000,
31'b0010000000000000000010100010000,
31'b0100001000000000110000000000100,
31'b1010000100100000001000000000000,
31'b1100000000000000010001100000000,
31'b0010010000000000000100000000011,
31'b1000101000000000010000000000100,
31'b0000010010000000000000000010100,
31'b0101000000000000000000010100000,
31'b0101000000000010000000010100000,
31'b0101000000000100000000010100000,
31'b1000110000010000000000000000001,
31'b1101100000000000000010000000000,
31'b0010010000001000000000000100100,
31'b1000000110000000000000100000000,
31'b1000110000001000000000000000001,
31'b0101000000010000000000010100000,
31'b0010010000000000000000000100100,
31'b1000110000000010000000000000001,
31'b1000110000000000000000000000001,
31'b0001000100010000000000011000000,
31'b1101000000000000100000001000000,
31'b0100000000001000100001000000010,
31'b0100000000000000010000000100100,
31'b0001000001000000100010000000000,
31'b1001101000000000000000010000000,
31'b0100000000000000100001000000010,
31'b0100000000001000010000000100100,
31'b0001000100000000000000011000000,
31'b0001001000000000000010000100000,
31'b1010100000000000001000010000000,
31'b0100001000000001100100000000000,
31'b0001000100001000000000011000000,
31'b0010010000100000000000000100100,
31'b1010010000000000000001100000000,
31'b1000110000100000000000000000001,
31'b1000000000000000000011000000100,
31'b1000000100000000001000000110000,
31'b1000000101010000000000100000000,
31'b0000010001000000000000000010100,
31'b0010000010000000000101000000000,
31'b0110000000010000000000010001000,
31'b0010000010000100000101000000000,
31'b0001110000100001000000000000000,
31'b1000000101000100000000100000000,
31'b0110000000001000000000010001000,
31'b1000000101000000000000100000000,
31'b1000010000100000001001000000000,
31'b0110000000000010000000010001000,
31'b0110000000000000000000010001000,
31'b1010000000000000000001010000001,
31'b1010000110000000001000000000000,
31'b0000010100000000000100000000000,
31'b0000010100000010000100000000000,
31'b0000010100000100000100000000000,
31'b0000000000000000000010100100000,
31'b0001000010000000100010000000000,
31'b0001110000000101000000000000000,
31'b0100100100000000100000100000000,
31'b0001110000000001000000000000000,
31'b0000010100010000000100000000000,
31'b1000010000000100001001000000000,
31'b1000010000000010001001000000000,
31'b1000010000000000001001000000000,
31'b0001010000000000001000001000010,
31'b1100000000000000001000001010000,
31'b1000100000000010000000110000000,
31'b1000100000000000000000110000000,
31'b1000000100010100000000100000000,
31'b0000010000000100000000000010100,
31'b1000000100010000000000100000000,
31'b0000010000000000000000000010100,
31'b0101000010000000000000010100000,
31'b0100000000000000000001001000100,
31'b1000000100011000000000100000000,
31'b0000101000000000000000101000000,
31'b1000000100000100000000100000000,
31'b1000010000000000000110000100000,
31'b1000000100000000000000100000000,
31'b1000000100000010000000100000000,
31'b1000000100001100000000100000000,
31'b0110000001000000000000010001000,
31'b1000000100001000000000100000000,
31'b1000110010000000000000000000001,
31'b0000010101000000000100000000000,
31'b0000010101000010000100000000000,
31'b1000000100110000000000100000000,
31'b0000010000100000000000000010100,
31'b0001010000000000010000010010000,
31'b1100000000000000010000010000010,
31'b1100000000000000000000101100000,
31'b0011001000000000000010000010000,
31'b0000000000000000001010000010000,
31'b0000000100000000000001000100100,
31'b1000000100100000000000100000000,
31'b1000010001000000001001000000000,
31'b0000000100000000110000000000010,
31'b0110000000000000010000000010100,
31'b1000000000000000001000000000011,
31'b1000100001000000000000110000000,
31'b1001010000000000000000000000000,
31'b0100000000000000000000000010010,
31'b0000000001000000000000001000001,
31'b0100000000000100000000000010010,
31'b0000000000000000000011000001000,
31'b0100000000001000000000000010010,
31'b0000000001001000000000001000001,
31'b1100000000000000000010000000001,
31'b0000000000000001000000110000000,
31'b0100000000010000000000000010010,
31'b0000000001010000000000001000001,
31'b0100100000000000000000010100001,
31'b0000000000010000000011000001000,
31'b0100000010000000000110010000000,
31'b0000000101000000000000100001100,
31'b1100000000010000000010000000001,
31'b0000001010000000000100000000000,
31'b0100000000100000000000000010010,
31'b0000001010000100000100000000000,
31'b0100001100000000100000000000001,
31'b0000001010001000000100000000000,
31'b0100001000000001000010100000000,
31'b0000101000000000000010000100001,
31'b1100000000100000000010000000001,
31'b0000001010010000000100000000000,
31'b0100001000000000000001010001000,
31'b1000001000000000000000010000001,
31'b1001000000000000001010000000100,
31'b0000001010011000000100000000000,
31'b0000000010000001000001000000010,
31'b1111000000000000010000000000000,
31'b0011000010000000001100000000000,
31'b0000000000000100000000001000001,
31'b0100000001000000000000000010010,
31'b0000000000000000000000001000001,
31'b0000000000000010000000001000001,
31'b0000000001000000000011000001000,
31'b1001000000000000000001000000011,
31'b0000000000001000000000001000001,
31'b1000010000000000000000000011000,
31'b0000000001000001000000110000000,
31'b0100000001010000000000000010010,
31'b0000000000010000000000001000001,
31'b0000100000000000010000100010000,
31'b0010000100000001000001000000001,
31'b0010001100000000000000000100100,
31'b0000000100000000000000100001100,
31'b1000101100000000000000000000001,
31'b0000001011000000000100000000000,
31'b0110001000000000000000001000100,
31'b0000000000100000000000001000001,
31'b0010000000000000100100000010000,
31'b0000001011001000000100000000000,
31'b0010100000000000100000010000100,
31'b0000000000101000000000001000001,
31'b1000010000100000000000000011000,
31'b0001000000000100000100100000000,
31'b0001010100000000000010000100000,
31'b0001000000000000000100100000000,
31'b0001000000000010000100100000000,
31'b0101110000000000100000000000000,
31'b0000100100000001000000100000000,
31'b0100000100000000000000000100001,
31'b0101000010000001000010000000000,
31'b0000001000100000000100000000000,
31'b0100000010000000000000000010010,
31'b0000001000100100000100000000000,
31'b0110000000000000000100000000101,
31'b0000001000101000000100000000000,
31'b0100000010001000000000000010010,
31'b0000101001000000010000000001000,
31'b1100000010000000000010000000001,
31'b0000001000110000000100000000000,
31'b0100000010010000000000000010010,
31'b1001000000100001000000001000000,
31'b0110000000001000000000000100010,
31'b0100001000000000000000100001010,
31'b0100000000000000000110010000000,
31'b0110000000000010000000000100010,
31'b0110000000000000000000000100010,
31'b0000001000000000000100000000000,
31'b0000001000000010000100000000000,
31'b0000001000000100000100000000000,
31'b0010000100000000000000001000010,
31'b0000001000001000000100000000000,
31'b0000001000001010000100000000000,
31'b0000100000000000001001001000000,
31'b0011000000010000001100000000000,
31'b0000001000010000000100000000000,
31'b0000001000010010000100000000000,
31'b1001000000000001000000001000000,
31'b1001000000000011000000001000000,
31'b0000001000011000000100000000000,
31'b0000000000000001000001000000010,
31'b1010101000000000000000000000010,
31'b0011000000000000001100000000000,
31'b0000001001100000000100000000000,
31'b0100000100000000100100001000000,
31'b0000000010000000000000001000001,
31'b0000001100000000000000000010100,
31'b0000101000000100010000000001000,
31'b0010100000000000010000100100000,
31'b0000101000000000010000000001000,
31'b1000010010000000000000000011000,
31'b1000000000000000000100011000000,
31'b1010010000000000000000000101000,
31'b1000011000000000000000100000000,
31'b1000011000000010000000100000000,
31'b1000010000000000101000000010000,
31'b0010000000000001001000010000000,
31'b1000100000000000000000001010100,
31'b0110000001000000000000000100010,
31'b0000001001000000000100000000000,
31'b0000001001000010000100000000000,
31'b0000001001000100000100000000000,
31'b0010000101000000000000001000010,
31'b0000001001001000000100000000000,
31'b0000001000000001010000000000100,
31'b0000101000100000010000000001000,
31'b1100000000000000010000000101000,
31'b0000010000000001000000000000001,
31'b0000010000000011000000000000001,
31'b0001000010000000000100100000000,
31'b0101000000001001000010000000000,
31'b0000010000001001000000000000001,
31'b0000000000000000100100000100000,
31'b0101000000000011000010000000000,
31'b0101000000000001000010000000000,
31'b0010000000000000100000000000100,
31'b0100000100000000000000000010010,
31'b0010000000000100100000000000100,
31'b0100001000100000100000000000001,
31'b0010000000001000100000000000100,
31'b0100000100001000000000000010010,
31'b0010000000001100100000000000100,
31'b1100000100000000000010000000001,
31'b0010000000010000100000000000100,
31'b0010010000000001000000000000010,
31'b0010000000010100100000000000100,
31'b0010010000000101000000000000010,
31'b0010000001000001000001000000001,
31'b0010010000001001000000000000010,
31'b0000000001000000000000100001100,
31'b1000101001000000000000000000001,
31'b0010000000100000100000000000100,
31'b0100001000000100100000000000001,
31'b0100001000000010100000000000001,
31'b0100001000000000100000000000001,
31'b1011000010000000000001000000000,
31'b0100000000000101010000000000010,
31'b0100000001010000000000000100001,
31'b0100000000000001010000000000010,
31'b0010100010000001001000000000000,
31'b0010100000000000000010001000100,
31'b1001000000000000000001000110000,
31'b1000001010000000001001000000000,
31'b0100100000000000011000001000000,
31'b0000100001000001000000100000000,
31'b0100000001000000000000000100001,
31'b0100000001000010000000000100001,
31'b0010000001000000100000000000100,
31'b0100000101000000000000000010010,
31'b0000000100000000000000001000001,
31'b0000001010000000000000000010100,
31'b0010000001001000100000000000100,
31'b0010001000010000000000000100100,
31'b0000000100001000000000001000001,
31'b1000101000010000000000000000001,
31'b0010000001010000100000000000100,
31'b0010010001000001000000000000010,
31'b0000000100010000000000001000001,
31'b1000101000001000000000000000001,
31'b0010000000000001000001000000001,
31'b0010001000000000000000000100100,
31'b0000000000000000000000100001100,
31'b1000101000000000000000000000001,
31'b0110000010000000000000000010001,
31'b1001000000000000001001100000000,
31'b0100000000000000000100000000110,
31'b0100001001000000100000000000001,
31'b0100100000000000000000010010010,
31'b0000100000010001000000100000000,
31'b0100000000010000000000000100001,
31'b0100000001000001010000000000010,
31'b0100100010000000000110000000000,
31'b0001010000000000000010000100000,
31'b0100000000001000000000000100001,
31'b0100010000000001100100000000000,
31'b0100000000000100000000000100001,
31'b0000100000000001000000100000000,
31'b0100000000000000000000000100001,
31'b0100000000000010000000000100001,
31'b0010000010000000100000000000100,
31'b0100000110000000000000000010010,
31'b0010000010000100100000000000100,
31'b0010000000100000000000001000010,
31'b1000000000000000100110000000000,
31'b1001100000000000000000100000001,
31'b1101000000000001000000000100000,
31'b0011000000000000000000100100100,
31'b0010100000100001001000000000000,
31'b0010010010000001000000000000010,
31'b0100100000000000001001000100000,
31'b0010000000000000001000000001100,
31'b1001000000000000010000001010000,
31'b1000100000100000000100001000000,
31'b0100000000000000010010000001000,
31'b0110000100000000000000000100010,
31'b0000001100000000000100000000000,
31'b0010000000000100000000001000010,
31'b0010000000000010000000001000010,
31'b0010000000000000000000001000010,
31'b1011000000000000000001000000000,
31'b1011000000000010000001000000000,
31'b1011000000000100000001000000000,
31'b0010000000001000000000001000010,
31'b0010100000000001001000000000000,
31'b1000100000001000000100001000000,
31'b1001000100000001000000001000000,
31'b1000001000000000001001000000000,
31'b1011000000010000000001000000000,
31'b1000100000000000000100001000000,
31'b0100000011000000000000000100001,
31'b1000100000000100000100001000000,
31'b0110000000100000000000000010001,
31'b0100000000000000100100001000000,
31'b0000001000000010000000000010100,
31'b0000001000000000000000000010100,
31'b1001000000000000001000010000010,
31'b0000101000000000000100010000000,
31'b0000110000000010000000101000000,
31'b0000110000000000000000101000000,
31'b1000010000000000010010000000010,
31'b1000001000000000000110000100000,
31'b1000011100000000000000100000000,
31'b1000000000000000010000001001000,
31'b0011000000000000001000000010100,
31'b0010001010000000000000000100100,
31'b0000010000000000010000000010001,
31'b1000101010000000000000000000001,
31'b0110000000000000000000000010001,
31'b0110000000000010000000000010001,
31'b0110000000000100000000000010001,
31'b0010000001000000000000001000010,
31'b1100000000000000000100010100000,
31'b0000101000100000000100010000000,
31'b1110000000000000000010000000010,
31'b0011010000000000000010000010000,
31'b0100100000000000000110000000000,
31'b0101000000000000100000100000001,
31'b0100100000000100000110000000000,
31'b1000001001000000001001000000000,
31'b0100100000001000000110000000000,
31'b0000100010000001000000100000000,
31'b0100000010000000000000000100001,
31'b0101000100000001000010000000000,
31'b0000000010100000000100000000000,
31'b0100001000000000000000000010010,
31'b0000001001000000000000001000001,
31'b0100001000000100000000000010010,
31'b0000001000000000000011000001000,
31'b0100001000001000000000000010010,
31'b0000100011000000010000000001000,
31'b1100001000000000000010000000001,
31'b0000001000000001000000110000000,
31'b0100001000010000000000000010010,
31'b1000000000100000000000010000001,
31'b1010010000001000001000000000000,
31'b0100000010000000000000100001010,
31'b1010010000000100001000000000000,
31'b1010010000000010001000000000000,
31'b1010010000000000001000000000000,
31'b0000000010000000000100000000000,
31'b0000000010000010000100000000000,
31'b0000000010000100000100000000000,
31'b0100000100000000100000000000001,
31'b0000000010001000000100000000000,
31'b0100000000000001000010100000000,
31'b0000100000000000000010000100001,
31'b0100000100001000100000000000001,
31'b0000000010010000000100000000000,
31'b0100000000000000000001010001000,
31'b1000000000000000000000010000001,
31'b1000000000000010000000010000001,
31'b0000000010011000000100000000000,
31'b0100000000010001000010100000000,
31'b1000000000001000000000010000001,
31'b1010010000100000001000000000000,
31'b0000001000000100000000001000001,
31'b0110000000100000000000001000100,
31'b0000001000000000000000001000001,
31'b0000001000000010000000001000001,
31'b0000100010000100010000000001000,
31'b0010000100010000000000000100100,
31'b0000100010000000010000000001000,
31'b1000100100010000000000000000001,
31'b1001000000000001000100000000001,
31'b0110000000000000001000000001010,
31'b1000010010000000000000100000000,
31'b1000100100001000000000000000001,
31'b0100100100000000000001000001000,
31'b0010000100000000000000000100100,
31'b1000100100000010000000000000001,
31'b1000100100000000000000000000001,
31'b0000000011000000000100000000000,
31'b0110000000000000000000001000100,
31'b0000001000100000000000001000001,
31'b0110000000000100000000001000100,
31'b0000000011001000000100000000000,
31'b0010000000000000001100100000000,
31'b0000100010100000010000000001000,
31'b0010010000000000000001000010100,
31'b0001010000000000000000011000000,
31'b0110000000010000000000001000100,
31'b1000000001000000000000010000001,
31'b1000100000000000001000100000010,
31'b0001010000001000000000011000000,
31'b0010000100100000000000000100100,
31'b1010000100000000000001100000000,
31'b1000100100100000000000000000001,
31'b0000000000100000000100000000000,
31'b0000000000100010000100000000000,
31'b0000000000100100000100000000000,
31'b0000000101000000000000000010100,
31'b0000000000101000000100000000000,
31'b0000000000101010000100000000000,
31'b0000100001000000010000000001000,
31'b0001100100100001000000000000000,
31'b0000000000110000000100000000000,
31'b0000000000110010000100000000000,
31'b1000010001000000000000100000000,
31'b1000010001000010000000100000000,
31'b0100000000000000000000100001010,
31'b0100001000000000000110010000000,
31'b1010100000100000000000000000010,
31'b1010010010000000001000000000000,
31'b0000000000000000000100000000000,
31'b0000000000000010000100000000000,
31'b0000000000000100000100000000000,
31'b0000000000000110000100000000000,
31'b0000000000001000000100000000000,
31'b0000000000001010000100000000000,
31'b0000000000001100000100000000000,
31'b0001100100000001000000000000000,
31'b0000000000010000000100000000000,
31'b0000000000010010000100000000000,
31'b0000000000010100000100000000000,
31'b1000000100000000001001000000000,
31'b0000000000011000000100000000000,
31'b0000001000000001000001000000010,
31'b1010100000000000000000000000010,
31'b1010100000000010000000000000010,
31'b0000000001100000000100000000000,
31'b0000000100000100000000000010100,
31'b0001000000000001000000010000000,
31'b0000000100000000000000000010100,
31'b0000100000000100010000000001000,
31'b0000100100000000000100010000000,
31'b0000100000000000010000000001000,
31'b0000100000000010010000000001000,
31'b1000010000000100000000100000000,
31'b1000010000000110000000100000000,
31'b1000010000000000000000100000000,
31'b1000010000000010000000100000000,
31'b1100100000000000100100000000000,
31'b0010001000000001001000010000000,
31'b1000010000001000000000100000000,
31'b1000100110000000000000000000001,
31'b0000000001000000000100000000000,
31'b0000000001000010000100000000000,
31'b0000000001000100000100000000000,
31'b0000000100100000000000000010100,
31'b0000000001001000000100000000000,
31'b0000000000000001010000000000100,
31'b0000100000100000010000000001000,
31'b0001000000000000000100000011000,
31'b0000000001010000000100000000000,
31'b0000010000000000000001000100100,
31'b1000010000100000000000100000000,
31'b1000010000100010000000100000000,
31'b0000010000000000110000000000010,
31'b0000001000000000100100000100000,
31'b1010100001000000000000000000010,
31'b0101001000000001000010000000000,
31'b0010001000000000100000000000100,
31'b0100001100000000000000000010010,
31'b0110000000000000000100001010000,
31'b0100000000100000100000000000001,
31'b0010010000000000000101000000000,
31'b0010010000000010000101000000000,
31'b0010010000000100000101000000000,
31'b1100000000000001001000000010000,
31'b0010001000010000100000000000100,
31'b0010011000000001000000000000010,
31'b1000110000000000000001000000010,
31'b1000100001001000000000000000001,
31'b0100100001000000000001000001000,
31'b0010000001000000000000000100100,
31'b1000100001000010000000000000001,
31'b1000100001000000000000000000001,
31'b0000000110000000000100000000000,
31'b0100000000000100100000000000001,
31'b0100000000000010100000000000001,
31'b0100000000000000100000000000001,
31'b0001010000000000100010000000000,
31'b0100000100000001000010100000000,
31'b0100010000000001000100000100000,
31'b0100000000001000100000000000001,
31'b0000000110010000000100000000000,
31'b1000000010000100001001000000000,
31'b1000000100000000000000010000001,
31'b1000000010000000001001000000000,
31'b0001010000010000100010000000000,
31'b0010010000000000000010100010000,
31'b1010000001000000000001100000000,
31'b1000100001100000000000000000001,
31'b0010001001000000100000000000100,
31'b0010000000000000000100000000011,
31'b0000001100000000000000001000001,
31'b0000000010000000000000000010100,
31'b0101010000000000000000010100000,
31'b0010000000010000000000000100100,
31'b1000100000010010000000000000001,
31'b1000100000010000000000000000001,
31'b0100100000001000000001000001000,
31'b0010000000001000000000000100100,
31'b1000100000001010000000000000001,
31'b1000100000001000000000000000001,
31'b0100100000000000000001000001000,
31'b0010000000000000000000000100100,
31'b1000100000000010000000000000001,
31'b1000100000000000000000000000001,
31'b0000000111000000000100000000000,
31'b0110000100000000000000001000100,
31'b0100001000000000000100000000110,
31'b0100000001000000100000000000001,
31'b0001010001000000100010000000000,
31'b0010000100000000001100100000000,
31'b1010000000010000000001100000000,
31'b1001000000000000100001000010000,
31'b0001010100000000000000011000000,
31'b0011000000000000000000101000010,
31'b1010000000001000000001100000000,
31'b1000100000101000000000000000001,
31'b1010000000000100000001100000000,
31'b0010000000100000000000000100100,
31'b1010000000000000000001100000000,
31'b1000100000100000000000000000001,
31'b0000000100100000000100000000000,
31'b0000000100100010000100000000000,
31'b0000000100100100000100000000000,
31'b0000000001000000000000000010100,
31'b0001000000000000000000000001100,
31'b0001000000000010000000000001100,
31'b0001000000000100000000000001100,
31'b0001100000100001000000000000000,
31'b0000000100110000000100000000000,
31'b1000000001000000000110000100000,
31'b1000010101000000000000100000000,
31'b1000000000100000001001000000000,
31'b0100000000000000000100001100000,
31'b0110010000000000000000010001000,
31'b0100001000000000010010000001000,
31'b1000100011000000000000000000001,
31'b0000000100000000000100000000000,
31'b0000000100000010000100000000000,
31'b0000000100000100000100000000000,
31'b0000000000000000010000010001000,
31'b0000000100001000000100000000000,
31'b0001100000000101000000000000000,
31'b0001100000000011000000000000000,
31'b0001100000000001000000000000000,
31'b0000000100010000000100000000000,
31'b1000000000000100001001000000000,
31'b1000000000000010001001000000000,
31'b1000000000000000001001000000000,
31'b0001000000000000001000001000010,
31'b1000101000000000000100001000000,
31'b1010100100000000000000000000010,
31'b1000000000001000001001000000000,
31'b0000000101100000000100000000000,
31'b0000000000000100000000000010100,
31'b0000000000000010000000000010100,
31'b0000000000000000000000000010100,
31'b0001000001000000000000000001100,
31'b0000100000000000000100010000000,
31'b0000100100000000010000000001000,
31'b0000000000001000000000000010100,
31'b1000010100000100000000100000000,
31'b1000000000000000000110000100000,
31'b1000010100000000000000100000000,
31'b0000000000010000000000000010100,
31'b0100100010000000000001000001000,
31'b0010000010000000000000000100100,
31'b1000100010000010000000000000001,
31'b1000100010000000000000000000001,
31'b0000000101000000000100000000000,
31'b0000000101000010000100000000000,
31'b0000000101000100000100000000000,
31'b0000000000100000000000000010100,
31'b0001000000000000010000010010000,
31'b0000100000100000000100010000000,
31'b0001100001000011000000000000000,
31'b0001100001000001000000000000000,
31'b0000010000000000001010000010000,
31'b1000000001000100001001000000000,
31'b1000010100100000000000100000000,
31'b1000000001000000001001000000000,
31'b0001000001000000001000001000010,
31'b0010000010100000000000000100100,
31'b1010000010000000000001100000000,
31'b1000100010100000000000000000001,
31'b1001100000000000000000000000000,
31'b1001100000000010000000000000000,
31'b1001100000000100000000000000000,
31'b1001100000000110000000000000000,
31'b1001100000001000000000000000000,
31'b1001100000001010000000000000000,
31'b1001100000001100000000000000000,
31'b1000000100000001000100000000000,
31'b1001100000010000000000000000000,
31'b1010000000000000000101001000000,
31'b1001100000010100000000000000000,
31'b0100010000000000000000010100001,
31'b0000000000000001001001000000000,
31'b0001001100000000000000001000000,
31'b0011000000000000000100000000010,
31'b1010101000000000001000000000000,
31'b1001100000100000000000000000000,
31'b1000000000000000010100000010000,
31'b1001100000100100000000000000000,
31'b1001000000000001000000000001100,
31'b1001100000101000000000000000000,
31'b1001000101000000000000010000000,
31'b0110000000010000001000000100000,
31'b1000100000000000010000010000100,
31'b1001100000110000000000000000000,
31'b1001000000000000100010001000000,
31'b0110000000001000001000000100000,
31'b0100000000000000100000000011000,
31'b0101000001000000100000000000000,
31'b0101000001000010100000000000000,
31'b0110000000000000001000000100000,
31'b0110000000000010001000000100000,
31'b1001100001000000000000000000000,
31'b1001100001000010000000000000000,
31'b1000000100000000010000000000100,
31'b1000100000001000000000000011000,
31'b1001100001001000000000000000000,
31'b1001000100100000000000010000000,
31'b1000100000000010000000000011000,
31'b1000100000000000000000000011000,
31'b1100000010000000000001000000100,
31'b0010000010000001000001100000000,
31'b1000101010000000000000100000000,
31'b0000010000000000010000100010000,
31'b0101000000100000100000000000000,
31'b0101000000100010100000000000000,
31'b0101000000100100100000000000000,
31'b1000100000010000000000000011000,
31'b1001100001100000000000000000000,
31'b1001000100001000000000010000000,
31'b1000100000000001000100010000000,
31'b0110001000000000101000000000000,
31'b1000000000000001000000000010100,
31'b1001000100000000000000010000000,
31'b1001000000000000010100000001000,
31'b1001000100000100000000010000000,
31'b0101000000001000100000000000000,
31'b0101000000001010100000000000000,
31'b0101000000001100100000000000000,
31'b0100000010000000000000100100000,
31'b0101000000000000100000000000000,
31'b0101000000000010100000000000000,
31'b0101000000000100100000000000000,
31'b0101000000000110100000000000000,
31'b1001100010000000000000000000000,
31'b1100010000000000000100000100000,
31'b1100000100000000000010100000000,
31'b0010000100000001000010000000100,
31'b1100000000000001100000000000001,
31'b0010000001000000000010010001000,
31'b0100001000100000100000100000000,
31'b0000000101000000000000101000000,
31'b1100000001000000000001000000100,
31'b0010000100000000100000001001000,
31'b1001000000000000000010000000110,
31'b0000000001000000000000000001101,
31'b0001000000000000000000000010101,
31'b0000000100000001000000010000001,
31'b0011000010000000000100000000010,
31'b0000000101010000000000101000000,
31'b0100000000000000001000000010000,
31'b0100000000000010001000000010000,
31'b0100000000000100001000000010000,
31'b0100000001010000000000100100000,
31'b0100000000001000001000000010000,
31'b0110000000000000100000000101000,
31'b0100001000000000100000100000000,
31'b0101000001000000001000000001000,
31'b0100000000010000001000000010000,
31'b0100000001000100000000100100000,
31'b0100000001000010000000100100000,
31'b0100000001000000000000100100000,
31'b0101000011000000100000000000000,
31'b1000010100000000000100001000000,
31'b1010011000000000000000000000010,
31'b1010000000000000010100000100000,
31'b1100000000010000000001000000100,
31'b0010000000010001000001100000000,
31'b1000101000010000000000100000000,
31'b0000000100001000000000101000000,
31'b0010001000000000000100100000010,
31'b0010000000000000000010010001000,
31'b0000011000000000010000000001000,
31'b0000000100000000000000101000000,
31'b1100000000000000000001000000100,
31'b0010000000000001000001100000000,
31'b1000101000000000000000100000000,
31'b0000000000000000000000000001101,
31'b1100000000001000000001000000100,
31'b0010000000010000000010010001000,
31'b1000101000001000000000100000000,
31'b0000000100010000000000101000000,
31'b0100000001000000001000000010000,
31'b0100000001000010001000000010000,
31'b0100000001000100001000000010000,
31'b0100000000010000000000100100000,
31'b1001000000000000001001000000001,
31'b1001000110000000000000010000000,
31'b0101000000000010001000000001000,
31'b0101000000000000001000000001000,
31'b0000100000000001000000000000001,
31'b0100000000000100000000100100000,
31'b0100000000000010000000100100000,
31'b0100000000000000000000100100000,
31'b0101000010000000100000000000000,
31'b0101000010000010100000000000000,
31'b0101000010000100100000000000000,
31'b0100000000001000000000100100000,
31'b1001100100000000000000000000000,
31'b1001100100000010000000000000000,
31'b0010000000000000001000001000000,
31'b1000000000001001000100000000000,
31'b1001100100001000000000000000000,
31'b1000000000000101000100000000000,
31'b1000000000000011000100000000000,
31'b1000000000000001000100000000000,
31'b1001100100010000000000000000000,
31'b0010100000000001000000000000010,
31'b1000001000000000000001000000010,
31'b1000001000000010000001000000010,
31'b0001001000000010000000001000000,
31'b0001001000000000000000001000000,
31'b1000001000001000000001000000010,
31'b1000000000010001000100000000000,
31'b1001100100100000000000000000000,
31'b1001000001001000000000010000000,
31'b1000000000000000000000010011000,
31'b1000000000101001000100000000000,
31'b1001000001000010000000010000000,
31'b1001000001000000000000010000000,
31'b1000000000100011000100000000000,
31'b1000000000100001000100000000000,
31'b0010010010000001001000000000000,
31'b0010100000100001000000000000010,
31'b0010000000000000000000000001110,
31'b0100100000000000000001000100010,
31'b0101000101000000100000000000000,
31'b0001001000100000000000001000000,
31'b0110000100000000001000000100000,
31'b1000001010000000000000110000000,
31'b1000000000000100010000000000100,
31'b1001000000101000000000010000000,
31'b1000000000000000010000000000100,
31'b1000000000000010010000000000100,
31'b1001000000100010000000010000000,
31'b1001000000100000000000010000000,
31'b1000000000001000010000000000100,
31'b0000000010000000000000101000000,
31'b1101001000000000000010000000000,
31'b0010100001000001000000000000010,
31'b1000000000010000010000000000100,
31'b1000011000001000000000000000001,
31'b0101000100100000100000000000000,
31'b0001001001000000000000001000000,
31'b1000011000000010000000000000001,
31'b1000011000000000000000000000001,
31'b1001000000001010000000010000000,
31'b1001000000001000000000010000000,
31'b1000000000100000010000000000100,
31'b1001000000001100000000010000000,
31'b1001000000000010000000010000000,
31'b1001000000000000000000010000000,
31'b1001000000000110000000010000000,
31'b1001000000000100000000010000000,
31'b0101000100001000100000000000000,
31'b0001100000000000000010000100000,
31'b1010001000000000001000010000000,
31'b0100100000000001100100000000000,
31'b0101000100000000100000000000000,
31'b0000010000000001000000100000000,
31'b0101000100000100100000000000000,
31'b0001000010000000000100000000001,
31'b1100000000000100000010100000000,
31'b0010000000010000100000001001000,
31'b1100000000000000000010100000000,
31'b0010000000000001000010000000100,
31'b0100000000000101011000000000000,
31'b0000000001000100000000101000000,
31'b0100000000000001011000000000000,
31'b0000000001000000000000101000000,
31'b0010010000100001001000000000000,
31'b0010000000000000100000001001000,
31'b1100000000010000000010100000000,
31'b0010000000010001000010000000100,
31'b0000000000000011000000010000001,
31'b0000000000000001000000010000001,
31'b0100100000000000000000110100000,
31'b0000000001010000000000101000000,
31'b0100000100000000001000000010000,
31'b0100000100000010001000000010000,
31'b1100000000100000000010100000000,
31'b0010110000000000000000001000010,
31'b0100000100001000001000000010000,
31'b1001000011000000000000010000000,
31'b0100001100000000100000100000000,
31'b0001011000000001000000000000000,
31'b0010010000000001001000000000000,
31'b1000010000001000000100001000000,
31'b0010010000000101001000000000000,
31'b1100000000000000000101000010000,
31'b1010000000000000000000010101000,
31'b1000010000000000000100001000000,
31'b1000001000000010000000110000000,
31'b1000001000000000000000110000000,
31'b1001000000000000000001100000010,
31'b0000000000001100000000101000000,
31'b1000000010000000010000000000100,
31'b0000000000001000000000101000000,
31'b0000000000000110000000101000000,
31'b0000000000000100000000101000000,
31'b0000000000000010000000101000000,
31'b0000000000000000000000101000000,
31'b1100000100000000000001000000100,
31'b0010000100000001000001100000000,
31'b1000101100000000000000100000000,
31'b0000000100000000000000000001101,
31'b0000100000000100010000000010001,
31'b0000000001000001000000010000001,
31'b0000100000000000010000000010001,
31'b0000000000010000000000101000000,
31'b0100010000010000000110000000000,
31'b1001000010001000000000010000000,
31'b1000000010100000010000000000100,
31'b0001000000000000000000000100110,
31'b1001000010000010000000010000000,
31'b1001000010000000000000010000000,
31'b0001000000000000110001000000000,
31'b0000000000100000000000101000000,
31'b0100010000000000000110000000000,
31'b0100010000000010000110000000000,
31'b0100010000000100000110000000000,
31'b0100000100000000000000100100000,
31'b0101000110000000100000000000000,
31'b0001000000000100000100000000001,
31'b0001000000000010000100000000001,
31'b0001000000000000000100000000001,
31'b1001101000000000000000000000000,
31'b0000000000000000001100000000010,
31'b1001101000000100000000000000000,
31'b0011000000000001000001000000000,
31'b1010000000000001000000001000010,
31'b0001000100010000000000001000000,
31'b0100000010100000100000100000000,
31'b1010100000010000001000000000000,
31'b1001101000010000000000000000000,
31'b0001000100001000000000001000000,
31'b1000000100000000000001000000010,
31'b1010100000001000001000000000000,
31'b0001000100000010000000001000000,
31'b0001000100000000000000001000000,
31'b1010100000000010001000000000000,
31'b1010100000000000001000000000000,
31'b0101000000000010000000000100000,
31'b0101000000000000000000000100000,
31'b0101000000000110000000000100000,
31'b0101000000000100000000000100000,
31'b0101000000001010000000000100000,
31'b0101000000001000000000000100000,
31'b0100000010000000100000100000000,
31'b0101000000001100000000000100000,
31'b0110000011000000000000000001000,
31'b0101000000010000000000000100000,
31'b1000110000000000000000010000001,
31'b0101000000010100000000000100000,
31'b0101001001000000100000000000000,
31'b0100000000000000001000100001000,
31'b1010010010000000000000000000010,
31'b1010100000100000001000000000000,
31'b1001101001000000000000000000000,
31'b0001000000000000100010010000000,
31'b1000100010010000000000100000000,
31'b0110000000100000101000000000000,
31'b0010000010000000000100100000010,
31'b0001000101010000000000001000000,
31'b0000010010000000010000000001000,
31'b1000101000000000000000000011000,
31'b1101000100000000000010000000000,
31'b0001000101001000000000001000000,
31'b1000100010000000000000100000000,
31'b1000100010000010000000100000000,
31'b0101001000100000100000000000000,
31'b0001000101000000000000001000000,
31'b1000100010001000000000100000000,
31'b1000010100000000000000000000001,
31'b0110000010010000000000000001000,
31'b0101000001000000000000000100000,
31'b0110000000000010101000000000000,
31'b0110000000000000101000000000000,
31'b1001000000000000000010001100000,
31'b1001001100000000000000010000000,
31'b0100000000000000000000000111000,
31'b0110000000001000101000000000000,
31'b0110000010000000000000000001000,
31'b0110000010000010000000000001000,
31'b1010000100000000001000010000000,
31'b1010000010000000000001000000001,
31'b0101001000000000100000000000000,
31'b0101001000000010100000000000000,
31'b0101001000000100100000000000000,
31'b1000100000000000000001010000010,
31'b1100000000000000010000000000010,
31'b0001010000000000010000000010000,
31'b1100000000000100010000000000010,
31'b0011000010000001000001000000000,
31'b1100000000001000010000000000010,
31'b0001010000001000010000000010000,
31'b0100000000100000100000100000000,
31'b0101000000000000010001001000000,
31'b1100000000010000010000000000010,
31'b0001010000010000010000000010000,
31'b1000100001000000000000100000000,
31'b1000100001000010000000100000000,
31'b0001001000000000000000000010101,
31'b0001000110000000000000001000000,
31'b1010010000100000000000000000010,
31'b1010100010000000001000000000000,
31'b0000110000000000000100000000000,
31'b0101000010000000000000000100000,
31'b0100000000001000100000100000000,
31'b0101000010000100000000000100000,
31'b0100000000000100100000100000000,
31'b0101000010001000000000000100000,
31'b0100000000000000100000100000000,
31'b0100000000000010100000100000000,
31'b0110000001000000000000000001000,
31'b0110000001000010000000000001000,
31'b1010010000001000000000000000010,
31'b1010000001000000000001000000001,
31'b1010010000000100000000000000010,
31'b1010000000000000000010001001000,
31'b1010010000000000000000000000010,
31'b1000000100000000000000110000000,
31'b1100000001000000010000000000010,
31'b0001010001000000010000000010000,
31'b1000100000010000000000100000000,
31'b1000100000010010000000100000000,
31'b0010000000000000000100100000010,
31'b0000010100000000000100010000000,
31'b0000010000000000010000000001000,
31'b0000010000000010010000000001000,
31'b1000100000000100000000100000000,
31'b1100000000000001000000000100001,
31'b1000100000000000000000100000000,
31'b1000100000000010000000100000000,
31'b1100010000000000100100000000000,
31'b0001000111000000000000001000000,
31'b1000100000001000000000100000000,
31'b1000100000001010000000100000000,
31'b0110000000010000000000000001000,
31'b0110000000010010000000000001000,
31'b1010000000000000110100000000000,
31'b1010000000010000000001000000001,
31'b0110000000011000000000000001000,
31'b1000000100000001000000001000001,
31'b0100000001000000100000100000000,
31'b0101001000000000001000000001000,
31'b0110000000000000000000000001000,
31'b0110000000000010000000000001000,
31'b1000100000100000000000100000000,
31'b1010000000000000000001000000001,
31'b0110000000001000000000000001000,
31'b0110000000001010000000000001000,
31'b1010010001000000000000000000010,
31'b1010000000001000000001000000001,
31'b1001101100000000000000000000000,
31'b0001000000011000000000001000000,
31'b1000000000010000000001000000010,
31'b1000001000001001000100000000000,
31'b0010100000000000000101000000000,
31'b0001000000010000000000001000000,
31'b1000001000000011000100000000000,
31'b1000001000000001000100000000000,
31'b1000000000000100000001000000010,
31'b0001000000001000000000001000000,
31'b1000000000000000000001000000010,
31'b1000000000000010000001000000010,
31'b0001000000000010000000001000000,
31'b0001000000000000000000001000000,
31'b1000000000001000000001000000010,
31'b0001000000000100000000001000000,
31'b0101000100000010000000000100000,
31'b0101000100000000000000000100000,
31'b1000001000000000000000010011000,
31'b0101000100000100000000000100000,
31'b0001100000000000100010000000000,
31'b0000000000000000000100100000001,
31'b0100100000000001000100000100000,
31'b0001010010000001000000000000000,
31'b1001000000000000100000010100000,
31'b0001000000101000000000001000000,
31'b1000000000100000000001000000010,
31'b1000000010001000000000110000000,
31'b0001000000100010000000001000000,
31'b0001000000100000000000001000000,
31'b1000000010000010000000110000000,
31'b1000000010000000000000110000000,
31'b1101000000010000000010000000000,
31'b0001000100000000100010010000000,
31'b1000001000000000010000000000100,
31'b1000010000011000000000000000001,
31'b0101100000000000000000010100000,
31'b0001000001010000000000001000000,
31'b1000010000010010000000000000001,
31'b1000010000010000000000000000001,
31'b1101000000000000000010000000000,
31'b0001000001001000000000001000000,
31'b0000000000000000000000001011000,
31'b1000010000001000000000000000001,
31'b0100010000000000000001000001000,
31'b0001000001000000000000001000000,
31'b1000010000000010000000000000001,
31'b1000010000000000000000000000001,
31'b0010000010000000001100000000001,
31'b1110000000000000010000000000001,
31'b0010000000000000010001000001000,
31'b0110000100000000101000000000000,
31'b1001001000000010000000010000000,
31'b1001001000000000000000010000000,
31'b0100100000000000100001000000010,
31'b1001001000000100000000010000000,
31'b1101000000100000000010000000000,
31'b0001101000000000000010000100000,
31'b1010000000000000001000010000000,
31'b1010000000000010001000010000000,
31'b0101001100000000100000000000000,
31'b0001000001100000000000001000000,
31'b1010000000001000001000010000000,
31'b1000010000100000000000000000001,
31'b1100000100000000010000000000010,
31'b0001010100000000010000000010000,
31'b1100001000000000000010100000000,
31'b0011000000000000000000001110000,
31'b0010100010000000000101000000000,
31'b0001000010010000000000001000000,
31'b0100001000000001011000000000000,
31'b0001010000100001000000000000000,
31'b1001000000000000010000100000100,
31'b0001000010001000000000001000000,
31'b1000000010000000000001000000010,
31'b1000000010000010000001000000010,
31'b0001000010000010000000001000000,
31'b0001000010000000000000001000000,
31'b1000000010001000000001000000010,
31'b1000000000100000000000110000000,
31'b0100000000000001000010000000001,
31'b0101000110000000000000000100000,
31'b0100000100001000100000100000000,
31'b0001010000001001000000000000000,
31'b0100000100000100100000100000000,
31'b0001010000000101000000000000000,
31'b0100000100000000100000100000000,
31'b0001010000000001000000000000000,
31'b0110000101000000000000000001000,
31'b1000000000001100000000110000000,
31'b1000000010100000000001000000010,
31'b1000000000001000000000110000000,
31'b1000000000000110000000110000000,
31'b1000000000000100000000110000000,
31'b1000000000000010000000110000000,
31'b1000000000000000000000110000000,
31'b0010000000100000001100000000001,
31'b0000010000001000000100010000000,
31'b1000100100010000000000100000000,
31'b0000110000000000000000000010100,
31'b0010000000000000000000001101000,
31'b0000010000000000000100010000000,
31'b0000010100000000010000000001000,
31'b0000001000000000000000101000000,
31'b1101000010000000000010000000000,
31'b0001000011001000000000001000000,
31'b1000100100000000000000100000000,
31'b1000100100000010000000100000000,
31'b0111000000000000000100000000100,
31'b0001000011000000000000001000000,
31'b1000100100001000000000100000000,
31'b1000010010000000000000000000001,
31'b0010000000000000001100000000001,
31'b1010000000000000100000010001000,
31'b0010000010000000010001000001000,
31'b0001010001001001000000000000000,
31'b1000000000000011000000001000001,
31'b1000000000000001000000001000001,
31'b0100000101000000100000100000000,
31'b0001010001000001000000000000000,
31'b0110000100000000000000000001000,
31'b0110000100000010000000000001000,
31'b1010000010000000001000010000000,
31'b1010000100000000000001000000001,
31'b0110000100001000000000000001000,
31'b1000000001000100000000110000000,
31'b1000100000000000001000000000011,
31'b1000000001000000000000110000000,
31'b0000000000000000011000000100000,
31'b0100100000000000000000000010010,
31'b0000100001000000000000001000001,
31'b0100100000000100000000000010010,
31'b0000100000000000000011000001000,
31'b0110000000000000000010000100100,
31'b0000100001001000000000001000001,
31'b1100100000000000000010000000001,
31'b0000100000000001000000110000000,
31'b0100100000010000000000000010010,
31'b0100000000000010000000010100001,
31'b0100000000000000000000010100001,
31'b0001000000000000010000100001000,
31'b0001011100000000000000001000000,
31'b0011010000000000000100000000010,
31'b1110000000000000000100000010000,
31'b0000101010000000000100000000000,
31'b1001000010000000001000000000010,
31'b0000101010000100000100000000000,
31'b0010000100000001100000000001000,
31'b0000101010001000000100000000000,
31'b0010000001000000100000010000100,
31'b0000001000000000000010000100001,
31'b0000000100000000000000011000001,
31'b0010001000000000000000010100100,
31'b0010000100000000000010001000100,
31'b1001000000000000100000000001010,
31'b0000000001000000100010000000001,
31'b0101010001000000100000000000000,
31'b0000000101000001000000100000000,
31'b1100000000000000100000001000001,
31'b0000000101000101000000100000000,
31'b0000100000000100000000001000001,
31'b0100100001000000000000000010010,
31'b0000100000000000000000001000001,
31'b0000100000000010000000001000001,
31'b0000100001000000000011000001000,
31'b0010000010000000010000100100000,
31'b0000100000001000000000001000001,
31'b1000110000000000000000000011000,
31'b0000100001000001000000110000000,
31'b0000000000000100010000100010000,
31'b0000100000010000000000001000001,
31'b0000000000000000010000100010000,
31'b0101010000100000100000000000000,
31'b0000001000000000111000000000000,
31'b1000001100000010000000000000001,
31'b1000001100000000000000000000001,
31'b0000101011000000000100000000000,
31'b0010000000001000100000010000100,
31'b0000100000100000000000001000001,
31'b0010000000000000000001101000000,
31'b1011000000000000000000100000010,
31'b0010000000000000100000010000100,
31'b0000100000101000000000001000001,
31'b0010000000001000000001101000000,
31'b0101010000001000100000000000000,
31'b0000000100001001000000100000000,
31'b0001100000000000000100100000000,
31'b0000000000000000100010000000001,
31'b0101010000000000100000000000000,
31'b0000000100000001000000100000000,
31'b0101010000000100100000000000000,
31'b0000000100000101000000100000000,
31'b0000101000100000000100000000000,
31'b1100000000000000000100000100000,
31'b0000101000100100000100000000000,
31'b1100000000000100000100000100000,
31'b0000101000101000000100000000000,
31'b1100000000001000000100000100000,
31'b0000001001000000010000000001000,
31'b0001001100100001000000000000000,
31'b0010001000000000110000100000000,
31'b1100000000010000000100000100000,
31'b0100000100000000001001000100000,
31'b0100000000000000000010000010100,
31'b0010000000000100011000000010000,
31'b1100000000000000000000000000111,
31'b0010000000000000011000000010000,
31'b0110100000000000000000000100010,
31'b0000101000000000000100000000000,
31'b1001000000000000001000000000010,
31'b0000101000000100000100000000000,
31'b1010000000000001000101000000000,
31'b0000101000001000000100000000000,
31'b1001000000001000001000000000010,
31'b0000000000000000001001001000000,
31'b0001001100000001000000000000000,
31'b0010000100000001001000000000000,
31'b1001000000010000001000000000010,
31'b1010001000001000000000000000010,
31'b0100010001000000000000100100000,
31'b1010001000000100000000000000010,
31'b1000000100000000000100001000000,
31'b1010001000000000000000000000010,
31'b1010001000000010000000000000010,
31'b0000101001100000000100000000000,
31'b1100000001000000000100000100000,
31'b0000100010000000000000001000001,
31'b0000101100000000000000000010100,
31'b0000001000000100010000000001000,
31'b0010000000000000010000100100000,
31'b0000001000000000010000000001000,
31'b0000010100000000000000101000000,
31'b1100010000000000000001000000100,
31'b0011000000000000011000000001000,
31'b1000111000000000000000100000000,
31'b0000010000000000000000000001101,
31'b1100001000000000100100000000000,
31'b0010100000000001001000010000000,
31'b1000000000000000000000001010100,
31'b1000001110000000000000000000001,
31'b0000101001000000000100000000000,
31'b1001000001000000001000000000010,
31'b0000101001000100000100000000000,
31'b1100000000000000001011000000000,
31'b0000101001001000000100000000000,
31'b0010000010000000100000010000100,
31'b0000001000100000010000000001000,
31'b0101010000000000001000000001000,
31'b0100000100000000000110000000000,
31'b0100010000000100000000100100000,
31'b0100010000000010000000100100000,
31'b0100010000000000000000100100000,
31'b0101010010000000100000000000000,
31'b0000100000000000100100000100000,
31'b1010001001000000000000000000010,
31'b0101100000000001000010000000000,
31'b0010100000000000100000000000100,
31'b0100100100000000000000000010010,
31'b1000000000000000100000000100001,
31'b1000010000001001000100000000000,
31'b0110000000000000001001000010000,
31'b1001000010000000000000100000001,
31'b1000010000000011000100000000000,
31'b1000010000000001000100000000000,
31'b0010100000010000100000000000100,
31'b0010110000000001000000000000010,
31'b1000011000000000000001000000010,
31'b1000001001001000000000000000001,
31'b0100001001000000000001000001000,
31'b0001011000000000000000001000000,
31'b1000001001000010000000000000001,
31'b1000001001000000000000000000001,
31'b0010100000100000100000000000100,
31'b0010000000010000000010001000100,
31'b1000010000000000000000010011000,
31'b0010000000000001100000000001000,
31'b0100000001000000000000010010010,
31'b0000000001010001000000100000000,
31'b0000000000000010000000011000001,
31'b0000000000000000000000011000001,
31'b0010000010000001001000000000000,
31'b0010000000000000000010001000100,
31'b0010010000000000000000000001110,
31'b0010000000010001100000000001000,
31'b0100000000000000011000001000000,
31'b0000000001000001000000100000000,
31'b0100100001000000000000000100001,
31'b0000000001000101000000100000000,
31'b1011000000000000001000000000001,
31'b0100000010000000000001100010000,
31'b1000010000000000010000000000100,
31'b1000010000000010010000000000100,
31'b0100001000010000000001000001000,
31'b0000001010000000000100010000000,
31'b1000010000001000010000000000100,
31'b1000001000010000000000000000001,
31'b0100001000001000000001000001000,
31'b0000001000000000000010000010010,
31'b1000010000010000010000000000100,
31'b1000001000001000000000000000001,
31'b0100001000000000000001000001000,
31'b0000000000100001000000100000000,
31'b1000001000000010000000000000001,
31'b1000001000000000000000000000001,
31'b0100000010010000000110000000000,
31'b0000000000011001000000100000000,
31'b1100000000000000000010010000001,
31'b0010000100000000000001101000000,
31'b0100000000000000000000010010010,
31'b0000000000010001000000100000000,
31'b0100100000010000000000000100001,
31'b0000000001000000000000011000001,
31'b0100000010000000000110000000000,
31'b0000000000001001000000100000000,
31'b0100100000001000000000000100001,
31'b0000000100000000100010000000001,
31'b0000000000000011000000100000000,
31'b0000000000000001000000100000000,
31'b0100100000000000000000000100001,
31'b0000000000000101000000100000000,
31'b0010100010000000100000000000100,
31'b1100000100000000000100000100000,
31'b1100010000000000000010100000000,
31'b0010100000100000000000001000010,
31'b1001000000000010000000100000001,
31'b1001000000000000000000100000001,
31'b0101000000000000000001100001000,
31'b0001001000100001000000000000000,
31'b0010000000100001001000000000000,
31'b1000000000101000000100001000000,
31'b0100000000000000001001000100000,
31'b0100000100000000000010000010100,
31'b1010000000000000100000000010001,
31'b1000000000100000000100001000000,
31'b0100100000000000010010000001000,
31'b1000001011000000000000000000001,
31'b0010000000010001001000000000000,
31'b1001000100000000001000000000010,
31'b0010100000000010000000001000010,
31'b0010100000000000000000001000010,
31'b1011100000000000000001000000000,
31'b1000000000010000000100001000000,
31'b0001001000000011000000000000000,
31'b0001001000000001000000000000000,
31'b0010000000000001001000000000000,
31'b1000000000001000000100001000000,
31'b0010000000000101001000000000000,
31'b1000101000000000001001000000000,
31'b1000000000000010000100001000000,
31'b1000000000000000000100001000000,
31'b1010001100000000000000000000010,
31'b1000000000000100000100001000000,
31'b0100000000110000000110000000000,
31'b0100000000000000000001100010000,
31'b1000010010000000010000000000100,
31'b0000101000000000000000000010100,
31'b0000001000000010000100010000000,
31'b0000001000000000000100010000000,
31'b0000010000000010000000101000000,
31'b0000010000000000000000101000000,
31'b0100000000100000000110000000000,
31'b0100000000100010000110000000000,
31'b0100000001000000001001000100000,
31'b1000100000000000010000001001000,
31'b0100001010000000000001000001000,
31'b0000001000010000000100010000000,
31'b1000001010000010000000000000001,
31'b1000001010000000000000000000001,
31'b0100000000010000000110000000000,
31'b0100000000100000000001100010000,
31'b1100000000000000000000000110100,
31'b0010100001000000000000001000010,
31'b0100000010000000000000010010010,
31'b0000001000100000000100010000000,
31'b0001010000000000110001000000000,
31'b0001001001000001000000000000000,
31'b0100000000000000000110000000000,
31'b0100000000000010000110000000000,
31'b0100000000000100000110000000000,
31'b0100010100000000000000100100000,
31'b0100000000001000000110000000000,
31'b0000000010000001000000100000000,
31'b0100100010000000000000000100001,
31'b0001010000000000000100000000001,
31'b0000100010100000000100000000000,
31'b0001000010000000010000000010000,
31'b0000101001000000000000001000001,
31'b0011010000000001000001000000000,
31'b0000101000000000000011000001000,
31'b0001010100010000000000001000000,
31'b0000000011000000010000000001000,
31'b1010000000000001000010000001000,
31'b0010000010000000110000100000000,
31'b0001010100001000000000001000000,
31'b1000100000100000000000010000001,
31'b1010000000000000000001110000000,
31'b0100000101000000000001000001000,
31'b0001010100000000000000001000000,
31'b1010000010100000000000000000010,
31'b1000000101000000000000000000001,
31'b0000100010000000000100000000000,
31'b0101010000000000000000000100000,
31'b0000100010000100000100000000000,
31'b0101010000000100000000000100000,
31'b0000100010001000000100000000000,
31'b0101010000001000000000000100000,
31'b0000000000000000000010000100001,
31'b0001000110000001000000000000000,
31'b0010000000000000000000010100100,
31'b0101010000010000000000000100000,
31'b1000100000000000000000010000001,
31'b1000100000000010000000010000001,
31'b1010000010000100000000000000010,
31'b0101000000000001010001000000000,
31'b1010000010000000000000000000010,
31'b1010000010000010000000000000010,
31'b0000101000000100000000001000001,
31'b0001010000000000100010010000000,
31'b0000101000000000000000001000001,
31'b1000000100011000000000000000001,
31'b0000000010000100010000000001000,
31'b0000000110000000000100010000000,
31'b0000000010000000010000000001000,
31'b1000000100010000000000000000001,
31'b0110000000000000100010000000100,
31'b0000000100000000000010000010010,
31'b1000110010000000000000100000000,
31'b1000000100001000000000000000001,
31'b0100000100000000000001000001000,
31'b0000000000000000111000000000000,
31'b1000000100000010000000000000001,
31'b1000000100000000000000000000001,
31'b0000100011000000000100000000000,
31'b0110100000000000000000001000100,
31'b0000101000100000000000001000001,
31'b1100000000000000000000001100001,
31'b0000100011001000000100000000000,
31'b0010100000000000001100100000000,
31'b0000000010100000010000000001000,
31'b1001000000000000000000000101010,
31'b0110010010000000000000000001000,
31'b1000000000000100001000100000010,
31'b1000100001000000000000010000001,
31'b1000000000000000001000100000010,
31'b0101011000000000100000000000000,
31'b0000001100000001000000100000000,
31'b1010000011000000000000000000010,
31'b1000000100100000000000000000001,
31'b0000100000100000000100000000000,
31'b0001000000000000010000000010000,
31'b0000100000100100000100000000000,
31'b0001000000000100010000000010000,
31'b0000100000101000000100000000000,
31'b0001000000001000010000000010000,
31'b0000000001000000010000000001000,
31'b0001000100100001000000000000000,
31'b0010000000000000110000100000000,
31'b0001000000010000010000000010000,
31'b1010000000101000000000000000010,
31'b0101000000000001000000001100000,
31'b1100000001000000100100000000000,
31'b0001010110000000000000001000000,
31'b1010000000100000000000000000010,
31'b1010000000100010000000000000010,
31'b0000100000000000000100000000000,
31'b0000100000000010000100000000000,
31'b0000100000000100000100000000000,
31'b0001000100001001000000000000000,
31'b0000100000001000000100000000000,
31'b0001000100000101000000000000000,
31'b0000000000000000000000010010100,
31'b0001000100000001000000000000000,
31'b0000100000010000000100000000000,
31'b0011000000000000000001001000000,
31'b1010000000001000000000000000010,
31'b1010000000001010000000000000010,
31'b1010000000000100000000000000010,
31'b1010000000000110000000000000010,
31'b1010000000000000000000000000010,
31'b1010000000000010000000000000010,
31'b0000100001100000000100000000000,
31'b0001000001000000010000000010000,
31'b0000000000001000010000000001000,
31'b0000100100000000000000000010100,
31'b0000000000000100010000000001000,
31'b0000000100000000000100010000000,
31'b0000000000000000010000000001000,
31'b0000000000000010010000000001000,
31'b1100000000001000100100000000000,
31'b0001000001010000010000000010000,
31'b1000110000000000000000100000000,
31'b1000110000000010000000100000000,
31'b1100000000000000100100000000000,
31'b0000000100010000000100010000000,
31'b0000000000010000010000000001000,
31'b1000000110000000000000000000001,
31'b0000100001000000000100000000000,
31'b0001000000000000000000010001100,
31'b0000100001000100000100000000000,
31'b0001000101001001000000000000000,
31'b0000100001001000000100000000000,
31'b0000100000000001010000000000100,
31'b0000000000100000010000000001000,
31'b0001000101000001000000000000000,
31'b0110010000000000000000000001000,
31'b0110010000000010000000000001000,
31'b1010000001001000000000000000010,
31'b1010010000000000000001000000001,
31'b1100000000100000100100000000000,
31'b0000101000000000100100000100000,
31'b1010000001000000000000000000010,
31'b1010000001000010000000000000010,
31'b0010101000000000100000000000100,
31'b0001010000011000000000001000000,
31'b1000010000010000000001000000010,
31'b1000000001011000000000000000001,
31'b0110000000000000000000011000100,
31'b0001010000010000000000001000000,
31'b1000000001010010000000000000001,
31'b1000000001010000000000000000001,
31'b1001000000000000000000000011001,
31'b0001010000001000000000001000000,
31'b1000010000000000000001000000010,
31'b1000000001001000000000000000001,
31'b0100000001000000000001000001000,
31'b0001010000000000000000001000000,
31'b1000000001000010000000000000001,
31'b1000000001000000000000000000001,
31'b0000100110000000000100000000000,
31'b0101010100000000000000000100000,
31'b0101000000000000000110100000000,
31'b0100100000000000100000000000001,
31'b0001110000000000100010000000000,
31'b0001000010000101000000000000000,
31'b0001000010000011000000000000000,
31'b0001000010000001000000000000000,
31'b0010001010000001001000000000000,
31'b0011000000000001000000000110000,
31'b1000100100000000000000010000001,
31'b1000100010000000001001000000000,
31'b0100001000000000011000001000000,
31'b0001010000100000000000001000000,
31'b1010000110000000000000000000010,
31'b1000000001100000000000000000001,
31'b0100000000011000000001000001000,
31'b0000000010001000000100010000000,
31'b1000011000000000010000000000100,
31'b1000000000011000000000000000001,
31'b0100000000010000000001000001000,
31'b0000000010000000000100010000000,
31'b1000000000010010000000000000001,
31'b1000000000010000000000000000001,
31'b0100000000001000000001000001000,
31'b0000000000000000000010000010010,
31'b1000000000001010000000000000001,
31'b1000000000001000000000000000001,
31'b0100000000000000000001000001000,
31'b1000000000000100000000000000001,
31'b1000000000000010000000000000001,
31'b1000000000000000000000000000001,
31'b0000000010000001000000000011000,
31'b0000001000011001000000100000000,
31'b0011000000000001001000100000000,
31'b1101000000000000001000000000100,
31'b0100001000000000000000010010010,
31'b0000001000010001000000100000000,
31'b1011000000000000010010000000000,
31'b1000000000110000000000000000001,
31'b0100001010000000000110000000000,
31'b0000001000001001000000100000000,
31'b1010010000000000001000010000000,
31'b1000000000101000000000000000001,
31'b0100000000100000000001000001000,
31'b0000001000000001000000100000000,
31'b1000000000100010000000000000001,
31'b1000000000100000000000000000001,
31'b0000100100100000000100000000000,
31'b0001000100000000010000000010000,
31'b0001000000101011000000000000000,
31'b0001000000101001000000000000000,
31'b0001100000000000000000000001100,
31'b0000000001000000000100010000000,
31'b0001000000100011000000000000000,
31'b0001000000100001000000000000000,
31'b0010001000100001001000000000000,
31'b0001010010001000000000001000000,
31'b1010000000000000001000100000001,
31'b1000100000100000001001000000000,
31'b0100100000000000000100001100000,
31'b0001010010000000000000001000000,
31'b1010000100100000000000000000010,
31'b1000000011000000000000000000001,
31'b0000100100000000000100000000000,
31'b0001000000001101000000000000000,
31'b0001000000001011000000000000000,
31'b0001000000001001000000000000000,
31'b0001000000000111000000000000000,
31'b0001000000000101000000000000000,
31'b0001000000000011000000000000000,
31'b0001000000000001000000000000000,
31'b0010001000000001001000000000000,
31'b1000100000000100001001000000000,
31'b1010000100001000000000000000010,
31'b1000100000000000001001000000000,
31'b1010000100000100000000000000010,
31'b1000001000000000000100001000000,
31'b1010000100000000000000000000010,
31'b0001000000010001000000000000000,
31'b0000000000100001000000000011000,
31'b0000000000001000000100010000000,
31'b0000100000000010000000000010100,
31'b0000100000000000000000000010100,
31'b0000000000000010000100010000000,
31'b0000000000000000000100010000000,
31'b0000000100000000010000000001000,
31'b0000000000000100000100010000000,
31'b0100001000100000000110000000000,
31'b0000000010000000000010000010010,
31'b1000110100000000000000100000000,
31'b1000000010001000000000000000001,
31'b0100000010000000000001000001000,
31'b0000000000010000000100010000000,
31'b1000000010000010000000000000001,
31'b1000000010000000000000000000001,
31'b0000000000000001000000000011000,
31'b0000000000101000000100010000000,
31'b0001000000000000010100000000100,
31'b0001000001001001000000000000000,
31'b0000000000100010000100010000000,
31'b0000000000100000000100010000000,
31'b0001000001000011000000000000000,
31'b0001000001000001000000000000000,
31'b0100001000000000000110000000000,
31'b0100001000000010000110000000000,
31'b0100001000000100000110000000000,
31'b1000100001000000001001000000000,
31'b0100001000001000000110000000000,
31'b0000001010000001000000100000000,
31'b1010000101000000000000000000010,
31'b1000000010100000000000000000001,
31'b1010000000000000000000000000000,
31'b1010000000000010000000000000000,
31'b1010000000000100000000000000000,
31'b1010000000000110000000000000000,
31'b1010000000001000000000000000000,
31'b1010000000001010000000000000000,
31'b1010000000001100000000000000000,
31'b1010000000001110000000000000000,
31'b1010000000010000000000000000000,
31'b1010000000010010000000000000000,
31'b1010000000010100000000000000000,
31'b1010000000010110000000000000000,
31'b1010000000011000000000000000000,
31'b1010000000011010000000000000000,
31'b0000100000000000000100000000010,
31'b1001001000000000001000000000000,
31'b1010000000100000000000000000000,
31'b1010000000100010000000000000000,
31'b1010000000100100000000000000000,
31'b1100001000000000000000000000101,
31'b1010000000101000000000000000000,
31'b1010000000101010000000000000000,
31'b1100010000010000010000000000000,
31'b0001000001000000001000011000000,
31'b1010000000110000000000000000000,
31'b1010000000110010000000000000000,
31'b1100010000001000010000000000000,
31'b0001000100000000101010000000000,
31'b1100010000000100010000000000000,
31'b0001000000000100010000000010010,
31'b1100010000000000010000000000000,
31'b0001000000000000010000000010010,
31'b1010000001000000000000000000000,
31'b1010000001000010000000000000000,
31'b1010000001000100000000000000000,
31'b1010000001000110000000000000000,
31'b1010000001001000000000000000000,
31'b1000000010000000001000100000000,
31'b1010000001001100000000000000000,
31'b1011000000000000000000000011000,
31'b1010000001010000000000000000000,
31'b1010000001010010000000000000000,
31'b1010000001010100000000000000000,
31'b0100000100000001000011000000000,
31'b1010000001011000000000000000000,
31'b1010001000000000100000000100000,
31'b1000000000000000100000100001000,
31'b1001001001000000001000000000000,
31'b1010000001100000000000000000000,
31'b1010000001100010000000000000000,
31'b1100000000000000100100000000010,
31'b0001010000000000100100000010000,
31'b1010000001101000000000000000000,
31'b1010100100000000000000010000000,
31'b0001000000000010001000011000000,
31'b0001000000000000001000011000000,
31'b0000000000000000010000000001010,
31'b0010000100000000000010000100000,
31'b0010010000000000000100100000000,
31'b0000010000000000010010001000000,
31'b0110100000000000100000000000000,
31'b0110100000000010100000000000000,
31'b1100010001000000010000000000000,
31'b0001000001000000010000000010010,
31'b1010000010000000000000000000000,
31'b1010000010000010000000000000000,
31'b1010000010000100000000000000000,
31'b1010000010000110000000000000000,
31'b0000000000000000000110000000100,
31'b1000000001000000001000100000000,
31'b1000000000010000000000000110000,
31'b1000000001000100001000100000000,
31'b1010000010010000000000000000000,
31'b1010000010010010000000000000000,
31'b1000000000001000000000000110000,
31'b1010000000000000101000000001000,
31'b1000000000000100000000000110000,
31'b1000000001010000001000100000000,
31'b1000000000000000000000000110000,
31'b1000000000000010000000000110000,
31'b1010000010100000000000000000000,
31'b1010000010100010000000000000000,
31'b1100000100000000000000001010000,
31'b0001010100000000000000001000010,
31'b1000010100000000000001000000000,
31'b1000010100000010000001000000000,
31'b1000010100000100000001000000000,
31'b0000010000010000001100000000000,
31'b1010000010110000000000000000000,
31'b0100100000000000101000100000000,
31'b1010010000000001000000001000000,
31'b0000010000001000001100000000000,
31'b1000010100010000000001000000000,
31'b0000010000000100001100000000000,
31'b1000000000100000000000000110000,
31'b0000010000000000001100000000000,
31'b1010000011000000000000000000000,
31'b0000000000000001010010000000000,
31'b1010000011000100000000000000000,
31'b1000001000000000100000000010000,
31'b1000000000000010001000100000000,
31'b1000000000000000001000100000000,
31'b1000000001010000000000000110000,
31'b1000000000000100001000100000000,
31'b1010000011010000000000000000000,
31'b1001000000000000000000000101000,
31'b1011001000000000000000100000000,
31'b1001000000000100000000000101000,
31'b1000000001000100000000000110000,
31'b1000000000010000001000100000000,
31'b1000000001000000000000000110000,
31'b1000000001000010000000000110000,
31'b1010000011100000000000000000000,
31'b1000000100000000000000000000011,
31'b0100100000000000100000000110000,
31'b0000000100001000000010000010000,
31'b1000010101000000000001000000000,
31'b1000000000100000001000100000000,
31'b0000000100000010000010000010000,
31'b0000000100000000000010000010000,
31'b0011000000000001000000000000001,
31'b1001000000100000000000000101000,
31'b0011000000000101000000000000001,
31'b0000010010000000010010001000000,
31'b0110100010000000100000000000000,
31'b1000000100000000000100000100100,
31'b1000010000000000000010100000100,
31'b0000010001000000001100000000000,
31'b1010000100000000000000000000000,
31'b1010000100000010000000000000000,
31'b1010000100000100000000000000000,
31'b1010000100000110000000000000000,
31'b1010000100001000000000000000000,
31'b1010000100001010000000000000000,
31'b1010000100001100000000000000000,
31'b0100000001000000000000110001000,
31'b1010000100010000000000000000000,
31'b0001000000000001000000000000010,
31'b1010000100010100000000000000000,
31'b0010000000000000001101000000000,
31'b1010000100011000000000000000000,
31'b0010101000000000000000001000000,
31'b1000000000000001000001001000000,
31'b1001001100000000001000000000000,
31'b1010000100100000000000000000000,
31'b1010000100100010000000000000000,
31'b1100000010000000000000001010000,
31'b0001010010000000000000001000010,
31'b1000010010000000000001000000000,
31'b1010100001000000000000010000000,
31'b1010000000000001010000000010000,
31'b0000010000000000110000010000000,
31'b1010000100110000000000000000000,
31'b0010000001000000000010000100000,
31'b0001100000000000000000000001110,
31'b0001000000000000101010000000000,
31'b1110000000000000000000001100000,
31'b0010101000100000000000001000000,
31'b1100010100000000010000000000000,
31'b0001000100000000010000000010010,
31'b1010000101000000000000000000000,
31'b1010000101000010000000000000000,
31'b1010000101000100000000000000000,
31'b0100000000010001000011000000000,
31'b1010000101001000000000000000000,
31'b1010100000100000000000010000000,
31'b0100001000000000000110000000010,
31'b0100000000000000000000110001000,
31'b1010000101010000000000000000000,
31'b0010000000100000000010000100000,
31'b0100001010000000000000010010000,
31'b0100000000000001000011000000000,
31'b0001010000000001000001000000001,
31'b0010101001000000000000001000000,
31'b0000000010000000000101100000000,
31'b0100000000010000000000110001000,
31'b1010000101100000000000000000000,
31'b1000000010000000000000000000011,
31'b0100000010000000000001000001010,
31'b0000000010001000000010000010000,
31'b1010100000000010000000010000000,
31'b1010100000000000000000010000000,
31'b0000001000000001000001010000000,
31'b0000000010000000000010000010000,
31'b0010000000000010000010000100000,
31'b0010000000000000000010000100000,
31'b0000001000000000000010100001000,
31'b0000000000000000000100010000010,
31'b0110100100000000100000000000000,
31'b0010000000001000000010000100000,
31'b0000001000010001000001010000000,
31'b0000000010010000000010000010000,
31'b1010000110000000000000000000000,
31'b1010000110000010000000000000000,
31'b1100000000100000000000001010000,
31'b0001100000000001000010000000100,
31'b1000010000100000000001000000000,
31'b1000010000100010000001000000000,
31'b1000010000100100000001000000000,
31'b0000010000000000000000100100100,
31'b1010000110010000000000000000000,
31'b0010000000000000010000000001001,
31'b1110000000000000010001000000000,
31'b0010000010000000001101000000000,
31'b1000010000110000000001000000000,
31'b0101001000000000000000010001000,
31'b1000000100000000000000000110000,
31'b1000000100000010000000000110000,
31'b0001000000000000000010000001000,
31'b1000000001000000000000000000011,
31'b1100000000000000000000001010000,
31'b0001010000000000000000001000010,
31'b1000010000000000000001000000000,
31'b1000010000000010000001000000000,
31'b1000010000000100000001000000000,
31'b0000000001000000000010000010000,
31'b1000000000000001010000000100000,
31'b1000000001010000000000000000011,
31'b1100000000010000000000001010000,
31'b0001010000010000000000001000010,
31'b1000010000010000000001000000000,
31'b1000010000010010000001000000000,
31'b1000010000010100000001000000000,
31'b0000010100000000001100000000000,
31'b1010000111000000000000000000000,
31'b1000000000100000000000000000011,
31'b0100001000010000000000010010000,
31'b0000001000000001000000100000010,
31'b1000010001100000000001000000000,
31'b1000000100000000001000100000000,
31'b0000000000100010000010000010000,
31'b0000000000100000000010000010000,
31'b0100110000000000100001000000000,
31'b1001000100000000000000000101000,
31'b0100001000000000000000010010000,
31'b0100001000000010000000010010000,
31'b0000010000000000001000000010100,
31'b1000000100010000001000100000000,
31'b0000000000000000000101100000000,
31'b0000000000110000000010000010000,
31'b1000000000000010000000000000011,
31'b1000000000000000000000000000011,
31'b0100000000000000000001000001010,
31'b0000000000001000000010000010000,
31'b1000010001000000000001000000000,
31'b0000000000000100000010000010000,
31'b0000000000000010000010000010000,
31'b0000000000000000000010000010000,
31'b1000000001000001010000000100000,
31'b1000000000010000000000000000011,
31'b0100001000100000000000010010000,
31'b0000000010000000000100010000010,
31'b1000010001010000000001000000000,
31'b1000000000000000000100000100100,
31'b0000000000100000000101100000000,
31'b0000000000010000000010000010000,
31'b1010001000000000000000000000000,
31'b1010001000000010000000000000000,
31'b1010001000000100000000000000000,
31'b0000100000000001000001000000000,
31'b1010001000001000000000000000000,
31'b1010001000001010000000000000000,
31'b1010001000001100000000000000000,
31'b1001000000010000001000000000000,
31'b1010001000010000000000000000000,
31'b1010001000010010000000000000000,
31'b1010001000010100000000000000000,
31'b1001000000001000001000000000000,
31'b1010001000011000000000000000000,
31'b1001000000000100001000000000000,
31'b1001000000000010001000000000000,
31'b1001000000000000001000000000000,
31'b0000000000000000000001000001100,
31'b0110100000000000000000000100000,
31'b0010000000000001000000100000001,
31'b1100000000000000000000000000101,
31'b0010000100000000100010000000000,
31'b0110100000001000000000000100000,
31'b0010000100000100100010000000000,
31'b1100000000001000000000000000101,
31'b0010000001000000000000011000000,
31'b0110100000010000000000000100000,
31'b0010000001000100000000011000000,
31'b1100000000010000000000000000101,
31'b0010000100010000100010000000000,
31'b1110000000000000000010010000000,
31'b1100011000000000010000000000000,
31'b1001000000100000001000000000000,
31'b1010001001000000000000000000000,
31'b1010001001000010000000000000000,
31'b1010001001000100000000000000000,
31'b1000000010000000100000000010000,
31'b1010001001001000000000000000000,
31'b1010000000010000100000000100000,
31'b0100010000000000010000011000000,
31'b1001000001010000001000000000000,
31'b1000000000000000001000000011000,
31'b1010000000001000100000000100000,
31'b1011000010000000000000100000000,
31'b1001000001001000001000000000000,
31'b1010000000000010100000000100000,
31'b1010000000000000100000000100000,
31'b1001000001000010001000000000000,
31'b1001000001000000001000000000000,
31'b0010000000010000000000011000000,
31'b0110100001000000000000000100000,
31'b0010000001000001000000100000001,
31'b1100000001000000000000000000101,
31'b0010000101000000100010000000000,
31'b0001010000000000001100100000000,
31'b0000000100000001000001010000000,
31'b0001000000000000000001000010100,
31'b0010000000000000000000011000000,
31'b0010000000000010000000011000000,
31'b0010000000000100000000011000000,
31'b0010000000000110000000011000000,
31'b0010000000001000000000011000000,
31'b1010000000100000100000000100000,
31'b0010000000001100000000011000000,
31'b1100000000000001100001000000000,
31'b1010001010000000000000000000000,
31'b1010001010000010000000000000000,
31'b1010001010000100000000000000000,
31'b1000000001000000100000000010000,
31'b1001000000000000100000000001000,
31'b1001000000000010100000000001000,
31'b1001000000000100100000000001000,
31'b1001000010010000001000000000000,
31'b1010001010010000000000000000000,
31'b0100100100000001010000000000000,
31'b1011000001000000000000100000000,
31'b1001000010001000001000000000000,
31'b1001000000010000100000000001000,
31'b1010000000000000000000100011000,
31'b1000001000000000000000000110000,
31'b1001000010000000001000000000000,
31'b0011010000000000000100000000000,
31'b0110100010000000000000000100000,
31'b0011010000000100000100000000000,
31'b1100000010000000000000000000101,
31'b1001000000100000100000000001000,
31'b0100100000010100000000000010000,
31'b0100100000010010000000000010000,
31'b0100100000010000000000000010000,
31'b0101100001000000000000000001000,
31'b0100000000000000000100010000100,
31'b0100100000001010000000000010000,
31'b0100100000001000000000000010000,
31'b0100100000000110000000000010000,
31'b0100100000000100000000000010000,
31'b0100100000000010000000000010000,
31'b0100100000000000000000000010000,
31'b1010001011000000000000000000000,
31'b1000000000000100100000000010000,
31'b1000000000000010100000000010000,
31'b1000000000000000100000000010000,
31'b1001000001000000100000000001000,
31'b1000001000000000001000100000000,
31'b1010000000000000001000000101000,
31'b1000000000001000100000000010000,
31'b1011000000000100000000100000000,
31'b1001001000000000000000000101000,
31'b1011000000000000000000100000000,
31'b1000000000010000100000000010000,
31'b0100100100000000000100000000100,
31'b1010000010000000100000000100000,
31'b1011000000001000000000100000000,
31'b1001000011000000001000000000000,
31'b0101100000010000000000000001000,
31'b1000001100000000000000000000011,
31'b1010000000000000000100001000001,
31'b1000000000100000100000000010000,
31'b0100100000000000001000100100000,
31'b0000000000000101001000000000001,
31'b0000000000000011001000000000001,
31'b0000000000000001001000000000001,
31'b0101100000000000000000000001000,
31'b0101100000000010000000000001000,
31'b1011000000100000000000100000000,
31'b1001100000000000000001000000001,
31'b0100000000000001010000010000000,
31'b0100100001000100000000000010000,
31'b0100100001000010000000000010000,
31'b0100100001000000000000000010000,
31'b1010001100000000000000000000000,
31'b1010001100000010000000000000000,
31'b1010001100000100000000000000000,
31'b1000000000000000000100001000010,
31'b0001000000000000000101000000000,
31'b0010100000010000000000001000000,
31'b0010000000000001001000000000010,
31'b1001000100010000001000000000000,
31'b1010001100010000000000000000000,
31'b0010100000001000000000001000000,
31'b0100010000000000110010000000000,
31'b1001000100001000001000000000000,
31'b0010100000000010000000001000000,
31'b0010100000000000000000001000000,
31'b1001000100000010001000000000000,
31'b1001000100000000001000000000000,
31'b0010000000001000100010000000000,
31'b0110100100000000000000000100000,
31'b0010000100000001000000100000001,
31'b1100000100000000000000000000101,
31'b0010000000000000100010000000000,
31'b0010000000000010100010000000000,
31'b0010000000000100100010000000000,
31'b0010110010000001000000000000000,
31'b0010000101000000000000011000000,
31'b0010100000101000000000001000000,
31'b0000000001000000000010100001000,
31'b1001000000000000000000100000011,
31'b0010000000010000100010000000000,
31'b0010100000100000000000001000000,
31'b0010000000010100100010000000000,
31'b1100000000000000000000101001000,
31'b1100000000000000000100000010001,
31'b0001010000000000000100000000011,
31'b0100000010010000000000010010000,
31'b0000000010000001000000100000010,
31'b0110000000000000000000010100000,
31'b0110000000000010000000010100000,
31'b0100000000000000000110000000010,
31'b0100001000000000000000110001000,
31'b1110100000000000000010000000000,
31'b0010100001001000000000001000000,
31'b0100000010000000000000010010000,
31'b0100001000000001000011000000000,
31'b0110000000010000000000010100000,
31'b0010100001000000000000001000000,
31'b0100000010001000000000010010000,
31'b1001000101000000001000000000000,
31'b0010000100010000000000011000000,
31'b1110000000000000100000001000000,
31'b0000000000010000000010100001000,
31'b0000001010001000000010000010000,
31'b0010000001000000100010000000000,
31'b1010101000000000000000010000000,
31'b0000000000000001000001010000000,
31'b0000001010000000000010000010000,
31'b0010000100000000000000011000000,
31'b0010001000000000000010000100000,
31'b0000000000000000000010100001000,
31'b0000001000000000000100010000010,
31'b0010000100001000000000011000000,
31'b0010100001100000000000001000000,
31'b0000000000010001000001010000000,
31'b0100000010000001000100000001000,
31'b1010001110000000000000000000000,
31'b0100100000010001010000000000000,
31'b0100000001010000000000010010000,
31'b0000100000000000000000001110000,
31'b0010010000000000000000000001100,
31'b0101000000010000000000010001000,
31'b0010010000000100000000000001100,
31'b0010110000100001000000000000000,
31'b0100100000000011010000000000000,
31'b0100100000000001010000000000000,
31'b0100000001000000000000010010000,
31'b0100100000000101010000000000000,
31'b0101000000000010000000010001000,
31'b0101000000000000000000010001000,
31'b1001000000000000000001010000001,
31'b1001000110000000001000000000000,
31'b1000000000000000100100000000100,
31'b1000001001000000000000000000011,
31'b1100001000000000000000001010000,
31'b0011000000000000000010100100000,
31'b1000011000000000000001000000000,
31'b1000011000000010000001000000000,
31'b1000100000000000100000010010000,
31'b0010110000000001000000000000000,
31'b1000001000000001010000000100000,
31'b1000010000000001000100000000010,
31'b0100000000000000010000000001100,
31'b0100100100001000000000000010000,
31'b1000011000010000000001000000000,
31'b0101000000100000000000010001000,
31'b0100100100000010000000000010000,
31'b0100100100000000000000000010000,
31'b0100100000000000000000000100011,
31'b0000000000000101000000100000010,
31'b0100000000010000000000010010000,
31'b0000000000000001000000100000010,
31'b0110000010000000000000010100000,
31'b1000001100000000001000100000000,
31'b0100000010000000000110000000010,
31'b0000001000100000000010000010000,
31'b0100000000000100000000010010000,
31'b0100100001000001010000000000000,
31'b0100000000000000000000010010000,
31'b0100000000000010000000010010000,
31'b0100100000000000000100000000100,
31'b0101000001000000000000010001000,
31'b0100000000001000000000010010000,
31'b0100000000100001000100000001000,
31'b1000001000000010000000000000011,
31'b1000001000000000000000000000011,
31'b0100001000000000000001000001010,
31'b0000001000001000000010000010000,
31'b1000011001000000000001000000000,
31'b1000000000000001110000000000000,
31'b0000001000000010000010000010000,
31'b0000001000000000000010000010000,
31'b0101100100000000000000000001000,
31'b1000010000000000100001000100000,
31'b0100000000100000000000010010000,
31'b0100000000100010000000010010000,
31'b1000010000000000010000000000110,
31'b1000001000000000000100000100100,
31'b0100000000101000000000010010000,
31'b0100000000000001000100000001000,
31'b1010010000000000000000000000000,
31'b1010010000000010000000000000000,
31'b1010010000000100000000000000000,
31'b1010010000000110000000000000000,
31'b1010010000001000000000000000000,
31'b1010010000001010000000000000000,
31'b1100000000110000010000000000000,
31'b0000101000010000010000000100000,
31'b1010010000010000000000000000000,
31'b1101000000000000000000010000100,
31'b1100000000101000010000000000000,
31'b0000101000001000010000000100000,
31'b1100000000100100010000000000000,
31'b0000101000000100010000000100000,
31'b1100000000100000010000000000000,
31'b0000101000000000010000000100000,
31'b1010010000100000000000000000000,
31'b1010010000100010000000000000000,
31'b1100000000011000010000000000000,
31'b0001000110000000000000001000010,
31'b0000000000000000100100000001000,
31'b1000000000000000001000010000001,
31'b1100000000010000010000000000000,
31'b0000000100000000110000010000000,
31'b1100000000001100010000000000000,
31'b0000101010000000000001001000000,
31'b1100000000001000010000000000000,
31'b0000000010001000001100000000000,
31'b1100000000000100010000000000000,
31'b0000000010000100001100000000000,
31'b1100000000000000010000000000000,
31'b0000000010000000001100000000000,
31'b1010010001000000000000000000000,
31'b1010010001000010000000000000000,
31'b0000100000000000110000000000000,
31'b0010000000000000000011000010000,
31'b1010010001001000000000000000000,
31'b1010000000000000000001000000011,
31'b0110000000000000000000000001010,
31'b0110000000000010000000000001010,
31'b1100100000000000000100000001000,
31'b0000100010000000011000000001000,
31'b0010000000100000000100100000000,
31'b0000100000000000000101000000001,
31'b0001000100000001000001000000001,
31'b0000001000000000001000001000001,
31'b1100000001100000010000000000000,
31'b0000101001000000010000000100000,
31'b1010010001100000000000000000000,
31'b0101001000000000000000001000100,
31'b0010000000010000000100100000000,
31'b0001000000000000100100000010000,
31'b1000100000000000000000100000010,
31'b1000100000000010000000100000010,
31'b1100000001010000010000000000000,
31'b0001010000000000001000011000000,
31'b0010000000000100000100100000000,
31'b0000001000000000000100000101000,
31'b0010000000000000000100100000000,
31'b0000000000000000010010001000000,
31'b1100000001000100010000000000000,
31'b0000001000100000001000001000001,
31'b1100000001000000010000000000000,
31'b0000000011000000001100000000000,
31'b1010010010000000000000000000000,
31'b1010010010000010000000000000000,
31'b1010010010000100000000000000000,
31'b0101000000000000000100000000101,
31'b1000000100100000000001000000000,
31'b1000010001000000001000100000000,
31'b1000010000010000000000000110000,
31'b0000000100000000000000100100100,
31'b1100000000000000000001001100000,
31'b0000101000100000000001001000000,
31'b1010000000100001000000001000000,
31'b0000000000101000001100000000000,
31'b1000010000000100000000000110000,
31'b0000000001000000000011000100000,
31'b1000010000000000000000000110000,
31'b0000000000100000001100000000000,
31'b1000000100001000000001000000000,
31'b1010100000000000001000000000010,
31'b1010000000010001000000001000000,
31'b0001000100000000000000001000010,
31'b1000000100000000000001000000000,
31'b1000000100000010000001000000000,
31'b1000000100000100000001000000000,
31'b0000000000010000001100000000000,
31'b1010000000000101000000001000000,
31'b0000101000000000000001001000000,
31'b1010000000000001000000001000000,
31'b0000000000001000001100000000000,
31'b1000000100010000000001000000000,
31'b0000000000000100001100000000000,
31'b0000000000000010001100000000000,
31'b0000000000000000001100000000000,
31'b1010010011000000000000000000000,
31'b1000100000000000000001010000000,
31'b0010001000000001000000010000000,
31'b1000100000000100000001010000000,
31'b1000010000000010001000100000000,
31'b1000010000000000001000100000000,
31'b0110000010000000000000000001010,
31'b1000010000000100001000100000000,
31'b0100100100000000100001000000000,
31'b0000100000000000011000000001000,
31'b0010001000010001000000010000000,
31'b0000100010000000000101000000001,
31'b0000000100000000001000000010100,
31'b0000000000000000000011000100000,
31'b1000010001000000000000000110000,
31'b0000000001100000001100000000000,
31'b1010000000000000000000110000001,
31'b1000100000100000000001010000000,
31'b0010001000100001000000010000000,
31'b0001000101000000000000001000010,
31'b1000000101000000000001000000000,
31'b1000010000100000001000100000000,
31'b1000000101000100000001000000000,
31'b0000010100000000000010000010000,
31'b0011010000000001000000000000001,
31'b0000101001000000000001001000000,
31'b0010000010000000000100100000000,
31'b0000000010000000010010001000000,
31'b1000000101010000000001000000000,
31'b0000000001000100001100000000000,
31'b1000000000000000000010100000100,
31'b0000000001000000001100000000000,
31'b0001000000000000100000000000100,
31'b1000000000000000000000110000010,
31'b1000000000000000010000001100000,
31'b1000000000000100000000110000010,
31'b1000000010100000000001000000000,
31'b1000000010100010000001000000000,
31'b1000000010100100000001000000000,
31'b0000000010000000000000100100100,
31'b1100000000000001000000000010000,
31'b0010000000000000000000100010100,
31'b1100000000000101000000000010000,
31'b0010010000000000001101000000000,
31'b1100000000001001000000000010000,
31'b0010111000000000000000001000000,
31'b1100000100100000010000000000000,
31'b0010100000000000000100110000000,
31'b1000000010001000000001000000000,
31'b1000000010001010000001000000000,
31'b1000000010001100000001000000000,
31'b0001000010000000000000001000010,
31'b1000000010000000000001000000000,
31'b1000000010000010000001000000000,
31'b1000000010000100000001000000000,
31'b0000000000000000110000010000000,
31'b1100000000100001000000000010000,
31'b0010010001000000000010000100000,
31'b1100000100001000010000000000000,
31'b0001010000000000101010000000000,
31'b1000000010010000000001000000000,
31'b1100000000000000000100010001000,
31'b1100000100000000010000000000000,
31'b0000000110000000001100000000000,
31'b1000100000000000001000000000001,
31'b1000100000000010001000000000001,
31'b0010000000000000001000000100100,
31'b0100100000000000001001000001000,
31'b1000100000001000001000000000001,
31'b0100001000000000000100001001000,
31'b0110000100000000000000000001010,
31'b0100000000000000010010000100000,
31'b1100000001000001000000000010000,
31'b0010010000100000000010000100000,
31'b0010000100100000000100100000000,
31'b1100100000000000010000010000000,
31'b0001000000000001000001000000001,
31'b0001001000000000000000000100100,
31'b0011000000000000000000100001100,
31'b1101000000000001000000000001000,
31'b1000100000100000001000000000001,
31'b1010000000000000001001100000000,
31'b0010000100010000000100100000000,
31'b0001000100000000100100000010000,
31'b1000000011000000000001000000000,
31'b1010110000000000000000010000000,
31'b1000101000000000010010000000000,
31'b0000010010000000000010000010000,
31'b0010010000000010000010000100000,
31'b0010010000000000000010000100000,
31'b0010000100000000000100100000000,
31'b0000010000000000000100010000010,
31'b1101100000000000000000000000100,
31'b0011100000000001000000100000000,
31'b1100000101000000010000000000000,
31'b0000010010010000000010000010000,
31'b1000000000101000000001000000000,
31'b1000000010000000000000110000010,
31'b1000000010000000010000001100000,
31'b0001000000100000000000001000010,
31'b1000000000100000000001000000000,
31'b1000000000100010000001000000000,
31'b1000000000100100000001000000000,
31'b0000000000000000000000100100100,
31'b1100000010000001000000000010000,
31'b0010010000000000010000000001001,
31'b0001100000000000100010000000010,
31'b0001000000000000001000000001100,
31'b1000000000110000000001000000000,
31'b1000000000110010000001000000000,
31'b1000010100000000000000000110000,
31'b0000000100100000001100000000000,
31'b1000000000001000000001000000000,
31'b1000000000001010000001000000000,
31'b1000000000001100000001000000000,
31'b0001000000000000000000001000010,
31'b1000000000000000000001000000000,
31'b1000000000000010000001000000000,
31'b1000000000000100000001000000000,
31'b0100000000000000000000000001001,
31'b1000000000011000000001000000000,
31'b1000001000000001000100000000010,
31'b1010000100000001000000001000000,
31'b0001000000010000000000001000010,
31'b1000000000010000000001000000000,
31'b1000000000010010000001000000000,
31'b1000000000010100000001000000000,
31'b0000000100000000001100000000000,
31'b1000100010000000001000000000001,
31'b1000100100000000000001010000000,
31'b0010001100000001000000010000000,
31'b0011001000000000000000000010100,
31'b1000000001100000000001000000000,
31'b1000010100000000001000100000000,
31'b1000000001100100000001000000000,
31'b0000010000100000000010000010000,
31'b0100100000000000100001000000000,
31'b0110000000000000010010000010000,
31'b0000100000000000001100010000000,
31'b1001001000000000000000010000010,
31'b0000000000000000001000000010100,
31'b0000000100000000000011000100000,
31'b0000010000000000000101100000000,
31'b0000010000110000000010000010000,
31'b1000000001001000000001000000000,
31'b1000010000000000000000000000011,
31'b1000000001001100000001000000000,
31'b0001000001000000000000001000010,
31'b1000000001000000000001000000000,
31'b1000000001000010000001000000000,
31'b1000000001000100000001000000000,
31'b0000010000000000000010000010000,
31'b1000000001011000000001000000000,
31'b1000010000010000000000000000011,
31'b0010100000000001100000000100000,
31'b0001000001010000000000001000010,
31'b1000000001010000000001000000000,
31'b1000010000000000000100000100100,
31'b1000000100000000000010100000100,
31'b0000010000010000000010000010000,
31'b1010011000000000000000000000000,
31'b1010011000000010000000000000000,
31'b1010011000000100000000000000000,
31'b1000000000000000010010010000000,
31'b1010011000001000000000000000000,
31'b0100100000000001000000001010000,
31'b0100000001000000010000011000000,
31'b0000100000010000010000000100000,
31'b1100000000000000001010000000001,
31'b0000100010100000000001001000000,
31'b0100000100000000110010000000000,
31'b0000100000001000010000000100000,
31'b0100000000000100001000000010010,
31'b0000100000000100010000000100000,
31'b0100000000000000001000000010010,
31'b0000100000000000010000000100000,
31'b0011000010000000000100000000000,
31'b0110110000000000000000000100000,
31'b0011000010000100000100000000000,
31'b1100010000000000000000000000101,
31'b1001000000000000000010000000100,
31'b1001000000000010000010000000100,
31'b1100001000010000010000000000000,
31'b0010100110000001000000000000000,
31'b0011000010010000000100000000000,
31'b0000100010000000000001001000000,
31'b1100001000001000010000000000000,
31'b0000100010000100000001001000000,
31'b1100001000000100010000000000000,
31'b0000100010001000000001001000000,
31'b1100001000000000010000000000000,
31'b0000100000100000010000000100000,
31'b1010011001000000000000000000000,
31'b0101000000100000000000001000100,
31'b0010000010000001000000010000000,
31'b1000010010000000100000000010000,
31'b0100000000000100010000011000000,
31'b0100000000000000000000100100010,
31'b0100000000000000010000011000000,
31'b0100000000000100000000100100010,
31'b1010000000000001000100000000001,
31'b0000000000100000000100000101000,
31'b0010001000100000000100100000000,
31'b0000101000000000000101000000001,
31'b0000000000000010001000001000001,
31'b0000000000000000001000001000001,
31'b0100000001000000001000000010010,
31'b0000100001000000010000000100000,
31'b0101000000000010000000001000100,
31'b0101000000000000000000001000100,
31'b0010001000010000000100100000000,
31'b1100000000000000110000000100000,
31'b1001000001000000000010000000100,
31'b0001000000000000001100100000000,
31'b1100000000000000000001000000110,
31'b0010000010000000000100000011000,
31'b0010010000000000000000011000000,
31'b0000000000000000000100000101000,
31'b0010001000000000000100100000000,
31'b0000001000000000010010001000000,
31'b0010010000001000000000011000000,
31'b0000000000100000001000001000001,
31'b1100001001000000010000000000000,
31'b0000100010000000000010000001001,
31'b0000000000000000100011000000000,
31'b0010100000000000010000000010000,
31'b0010000001000001000000010000000,
31'b1000010001000000100000000010000,
31'b0010000100000000000000000001100,
31'b0100100100000000000001000100000,
31'b0010000100000100000000000001100,
31'b0010100100100001000000000000000,
31'b0010000000000000000000101000001,
31'b0000100000100000000001001000000,
31'b0010000001010001000000010000000,
31'b0000100010001000010000000100000,
31'b0010000100010000000000000001100,
31'b0000100010000100010000000100000,
31'b1001100000100000000000000000010,
31'b0000100010000000010000000100000,
31'b0011000000000000000100000000000,
31'b0011000000000010000100000000000,
31'b0011000000000100000100000000000,
31'b0011000000000110000100000000000,
31'b1000001100000000000001000000000,
31'b1001000000000001001000001000000,
31'b1001100000010000000000000000010,
31'b0010100100000001000000000000000,
31'b0011000000010000000100000000000,
31'b0000100000000000000001001000000,
31'b1010001000000001000000001000000,
31'b0000100000000100000001001000000,
31'b1001100000000100000000000000010,
31'b0000100000001000000001001000000,
31'b1001100000000000000000000000010,
31'b0000001000000000001100000000000,
31'b0010000000000101000000010000000,
31'b1000101000000000000001010000000,
31'b0010000000000001000000010000000,
31'b1000010000000000100000000010000,
31'b0010000101000000000000000001100,
31'b1100000000000000100001001000000,
31'b0010000000001001000000010000000,
31'b1000010000001000100000000010000,
31'b0010000001000000000000101000001,
31'b0000101000000000011000000001000,
31'b0010000000010001000000010000000,
31'b1001000100000000000000010000010,
31'b0000000100000000000001011000000,
31'b0000001000000000000011000100000,
31'b0010000000011001000000010000000,
31'b0000100011000000010000000100000,
31'b0100000000000000000001010100000,
31'b0101000010000000000000001000100,
31'b0010000000100001000000010000000,
31'b1000010000100000100000000010000,
31'b1101000000000000010000100000000,
31'b0011000000000001010000000000100,
31'b0010000000101001000000010000000,
31'b0010000000000000000100000011000,
31'b0101110000000000000000000001000,
31'b0000100001000000000001001000000,
31'b0010001010000000000100100000000,
31'b0000100001000100000001001000000,
31'b1100100000000000000011000000000,
31'b0000100001001000000001001000000,
31'b1001100001000000000000000000010,
31'b0000100000000000000010000001001,
31'b1000000000000000000110000001000,
31'b1000001000000000000000110000010,
31'b1000001000000000010000001100000,
31'b1000010000000000000100001000010,
31'b0010000010000000000000000001100,
31'b0100100010000000000001000100000,
31'b0010010000000001001000000000010,
31'b0010100010100001000000000000000,
31'b1100001000000001000000000010000,
31'b0010110000001000000000001000000,
31'b0100000000000000110010000000000,
31'b0110100000000000000001000010000,
31'b0010110000000010000000001000000,
31'b0010110000000000000000001000000,
31'b0100000100000000001000000010010,
31'b0010000000000000101000000000100,
31'b1000001010001000000001000000000,
31'b0100100000000100010000001000000,
31'b0100100000000010010000001000000,
31'b0100100000000000010000001000000,
31'b1000001010000000000001000000000,
31'b1000001010000010000001000000000,
31'b1000100001000000010010000000000,
31'b0010100010000001000000000000000,
31'b0100000000000100000000100010001,
31'b0000100000000001000000000110000,
31'b0100000000000000000000100010001,
31'b0100100000010000010000001000000,
31'b1100000000000000000010100000010,
31'b0010110000100000000000001000000,
31'b1100001100000000010000000000000,
31'b0010100010010001000000000000000,
31'b1000101000000000001000000000001,
31'b0001000000000000000100000000011,
31'b0010001000000000001000000100100,
31'b0011000010000000000000000010100,
31'b0110010000000000000000010100000,
31'b0100000000000000000100001001000,
31'b1000100000100000010010000000000,
31'b1001000000000000000110000010000,
31'b0001000000001010000000000100100,
31'b0001000000001000000000000100100,
31'b0000000010000000100000100000100,
31'b1001000010000000000000010000010,
31'b0001000000000010000000000100100,
31'b0001000000000000000000000100100,
31'b1001000000100000000001100000000,
31'b1000000000000000110000001000000,
31'b0100000000000010001000000100001,
31'b0100000000000000001000000100001,
31'b0000100000000001001000100000000,
31'b0100100001000000010000001000000,
31'b1000100000000100010010000000000,
31'b0100000000100000000100001001000,
31'b1000100000000000010010000000000,
31'b1010000000000000100001000010000,
31'b0000000000000100010000010100000,
31'b0000000000000000000000101000010,
31'b0000000000000000010000010100000,
31'b0000000000000100000000101000010,
31'b1001000000000100000001100000000,
31'b0001000000100000000000000100100,
31'b1001000000000000000001100000000,
31'b1001000000000010000001100000000,
31'b0010000000001000000000000001100,
31'b0100100000001000000001000100000,
31'b0010000101000001000000010000000,
31'b0011000001000000000000000010100,
31'b0010000000000000000000000001100,
31'b0100100000000000000001000100000,
31'b0010000000000100000000000001100,
31'b0010100000100001000000000000000,
31'b0010000100000000000000101000001,
31'b1100000000000000000011010000000,
31'b0000000001000000100000100000100,
31'b1001000001000000000000010000010,
31'b0010000000010000000000000001100,
31'b0101010000000000000000010001000,
31'b0010000000010100000000000001100,
31'b0010100000110001000000000000000,
31'b1000001000001000000001000000000,
31'b1000001000001010000001000000000,
31'b1000100000000000001100001000000,
31'b0010100000001001000000000000000,
31'b1000001000000000000001000000000,
31'b1000001000000010000001000000000,
31'b1000001000000100000001000000000,
31'b0010100000000001000000000000000,
31'b1000001000011000000001000000000,
31'b1000000000000001000100000000010,
31'b0100010000000000010000000001100,
31'b1011000000000000001001000000000,
31'b1000001000010000000001000000000,
31'b1000001000010010000001000000000,
31'b1001100100000000000000000000010,
31'b0010100000010001000000000000000,
31'b0010000100000101000000010000000,
31'b0011000000000100000000000010100,
31'b0010000100000001000000010000000,
31'b0011000000000000000000000010100,
31'b0010000001000000000000000001100,
31'b0100100001000000000001000100000,
31'b0010000100001001000000010000000,
31'b0011000000001000000000000010100,
31'b0000000000001000000001011000000,
31'b1001000000000100000000010000010,
31'b0000000000000000100000100000100,
31'b1001000000000000000000010000010,
31'b0000000000000000000001011000000,
31'b0001000010000000000000000100100,
31'b0000000000001000100000100000100,
31'b1001000000001000000000010000010,
31'b1000001001001000000001000000000,
31'b1000011000000000000000000000011,
31'b0010100000000000010100000000100,
31'b0011000000100000000000000010100,
31'b1000001001000000000001000000000,
31'b1000010000000001110000000000000,
31'b1000100010000000010010000000000,
31'b0010100001000001000000000000000,
31'b1000000000001000010000000000110,
31'b1000000000000000100001000100000,
31'b0000000010000000010000010100000,
31'b1001000000100000000000010000010,
31'b1000000000000000010000000000110,
31'b1000000000001000100001000100000,
31'b1001000010000000000001100000000,
31'b0110000000000000001000000010001,
31'b1010100000000000000000000000000,
31'b1010100000000010000000000000000,
31'b0000000000000000000000000100101,
31'b0000001000000001000001000000000,
31'b1010100000001000000000000000000,
31'b1010100000001010000000000000000,
31'b0000000000010000000100000000010,
31'b0000001000001001000001000000000,
31'b1010100000010000000000000000000,
31'b1010100000010010000000000000000,
31'b0000000000001000000100000000010,
31'b0000001000010001000001000000000,
31'b0000000000000100000100000000010,
31'b0010001100000000000000001000000,
31'b0000000000000000000100000000010,
31'b0000000000000010000100000000010,
31'b1010100000100000000000000000000,
31'b1000000000000000000001100000001,
31'b0100000000000000000000100001000,
31'b0100000000000010000000100001000,
31'b1010100000101000000000000000000,
31'b1010000101000000000000010000000,
31'b0100000000001000000000100001000,
31'b0100001010010000000000000010000,
31'b1010100000110000000000000000000,
31'b1010000000000000100010001000000,
31'b0100000000010000000000100001000,
31'b0100001010001000000000000010000,
31'b0110000001000000100000000000000,
31'b0110000001000010100000000000000,
31'b0000000000100000000100000000010,
31'b0100001010000000000000000010000,
31'b1010100001000000000000000000000,
31'b1010100001000010000000000000000,
31'b0000010000000000110000000000000,
31'b0000010000000010110000000000000,
31'b1010100001001000000000000000000,
31'b1010000100100000000000010000000,
31'b0000010000001000110000000000000,
31'b0000010000001010110000000000000,
31'b1100010000000000000100000001000,
31'b0001000010000001000001100000000,
31'b0000010000010000110000000000000,
31'b0000010000000000000101000000001,
31'b0110000000100000100000000000000,
31'b0110000000100010100000000000000,
31'b0000000001000000000100000000010,
31'b0000001000000000100000000000101,
31'b1010100001100000000000000000000,
31'b1010000100001000000000010000000,
31'b0100000001000000000000100001000,
31'b0101001000000000101000000000000,
31'b1000010000000000000000100000010,
31'b1010000100000000000000010000000,
31'b1010000000000000010100000001000,
31'b1010000100000100000000010000000,
31'b0110000000001000100000000000000,
31'b0110000000001010100000000000000,
31'b0110000000001100100000000000000,
31'b1000000100000000000010000000101,
31'b0110000000000000100000000000000,
31'b0110000000000010100000000000000,
31'b0110000000000100100000000000000,
31'b0110000000000110100000000000000,
31'b1010100010000000000000000000000,
31'b1010100010000010000000000000000,
31'b0000000000000000000010010010000,
31'b0000001010000001000001000000000,
31'b1000000000000000000000010000011,
31'b1000100001000000001000100000000,
31'b0000000010010000000100000000010,
31'b0100001000110000000000000010000,
31'b1010100010010000000000000000000,
31'b0100001100000001010000000000000,
31'b0000000010001000000100000000010,
31'b0100001000101000000000000010000,
31'b0010000000000000000000000010101,
31'b0100001000100100000000000010000,
31'b0000000010000000000100000000010,
31'b0100001000100000000000000010000,
31'b1010100010100000000000000000000,
31'b1010010000000000001000000000010,
31'b0100000010000000000000100001000,
31'b0100001000011000000000000010000,
31'b1000110100000000000001000000000,
31'b0101000000000000100000000101000,
31'b0100001000010010000000000010000,
31'b0100001000010000000000000010000,
31'b0101001001000000000000000001000,
31'b0100000000000000101000100000000,
31'b0100001000001010000000000010000,
31'b0100001000001000000000000010000,
31'b0110000011000000100000000000000,
31'b0100001000000100000000000010000,
31'b0100001000000010000000000010000,
31'b0100001000000000000000000010000,
31'b1010100011000000000000000000000,
31'b1000010000000000000001010000000,
31'b0000010010000000110000000000000,
31'b1000101000000000100000000010000,
31'b1000100000000010001000100000000,
31'b1000100000000000001000100000000,
31'b0001010000000000000000011000010,
31'b1100000000000000000000011010000,
31'b0101001000100000000000000001000,
31'b0001000000000001000001100000000,
31'b0000010100000000001100010000000,
31'b0011000000000000000000000001101,
31'b0110000010100000100000000000000,
31'b1000100000010000001000100000000,
31'b0000000100000000100000001010000,
31'b0110000000000000000000001000110,
31'b0101001000010000000000000001000,
31'b1000100100000000000000000000011,
31'b0100000000000000100000000110000,
31'b0110000000001000001000000001000,
31'b1010000000000000001001000000001,
31'b1010000110000000000000010000000,
31'b0110000000000010001000000001000,
31'b0110000000000000001000000001000,
31'b0101001000000000000000000001000,
31'b0101001000000010000000000001000,
31'b1001000000000001000000000100100,
31'b1001001000000000000001000000001,
31'b0110000010000000100000000000000,
31'b0110000010000010100000000000000,
31'b0110000010000100100000000000000,
31'b0100001001000000000000000010000,
31'b1010100100000000000000000000000,
31'b1010100100000010000000000000000,
31'b0001000000000000001000001000000,
31'b0001000000000010001000001000000,
31'b1010100100001000000000000000000,
31'b1000000000000000001001000000010,
31'b0001000000001000001000001000000,
31'b1011000000000001000100000000000,
31'b1010100100010000000000000000000,
31'b0010001000001000000000001000000,
31'b0001000000010000001000001000000,
31'b0010100000000000001101000000000,
31'b0010001000000010000000001000000,
31'b0010001000000000000000001000000,
31'b0000000100000000000100000000010,
31'b0010001000000100000000001000000,
31'b1010100100100000000000000000000,
31'b1010000001001000000000010000000,
31'b0100000100000000000000100001000,
31'b0100011000000000010000001000000,
31'b1010000001000010000000010000000,
31'b1010000001000000000000010000000,
31'b0100000100001000000000100001000,
31'b1010000001000100000000010000000,
31'b0001010010000001001000000000000,
31'b0010100001000000000010000100000,
31'b0001000000000000000000000001110,
31'b1000000001000000000010000000101,
31'b0110000101000000100000000000000,
31'b0010001000100000000000001000000,
31'b0100000000000000000000001000101,
31'b0100001110000000000000000010000,
31'b1000010000000000001000000000001,
31'b1010000000101000000000010000000,
31'b0001000001000000001000001000000,
31'b0101000000000001010000100000000,
31'b1010000000100010000000010000000,
31'b1010000000100000000000010000000,
31'b0001000010000000010110000000000,
31'b1101000000000000001010000000000,
31'b1110001000000000000010000000000,
31'b0010100000100000000010000100000,
31'b0001000001010000001000001000000,
31'b1100010000000000010000010000000,
31'b0110000100100000100000000000000,
31'b0010001001000000000000001000000,
31'b0000000101000000000100000000010,
31'b0010001001000100000000001000000,
31'b1010000000001010000000010000000,
31'b1010000000001000000000010000000,
31'b0100000101000000000000100001000,
31'b1010000000001100000000010000000,
31'b1010000000000010000000010000000,
31'b1010000000000000000000010000000,
31'b1010000000000110000000010000000,
31'b1010000000000100000000010000000,
31'b0110000100001000100000000000000,
31'b0010100000000000000010000100000,
31'b1001001000000000001000010000000,
31'b1000000000000000000010000000101,
31'b0110000100000000100000000000000,
31'b0000000000000000000000000010110,
31'b0110000100000100100000000000000,
31'b0010000010000000000100000000001,
31'b1010100110000000000000000000000,
31'b0100001000010001010000000000000,
31'b0001000010000000001000001000000,
31'b0001000000000001000010000000100,
31'b1000110000100000000001000000000,
31'b1010010000000000000000100000001,
31'b0001000010001000001000001000000,
31'b0011000001000000000000101000000,
31'b0100010001000000100001000000000,
31'b0100001000000001010000000000000,
31'b0001010000000000100010000000010,
31'b1100000000000000100010000010000,
31'b0100001001000000000100000000100,
31'b0100000000000000100000000000011,
31'b0000000110000000000100000000010,
31'b0100001100100000000000000010000,
31'b1000000000000000001000110000000,
31'b1000100001000000000000000000011,
31'b1100100000000000000000001010000,
31'b0010011000001001000000000000000,
31'b1000110000000000000001000000000,
31'b1010000011000000000000010000000,
31'b1000110000000100000001000000000,
31'b0010011000000001000000000000000,
31'b0001010000000001001000000000000,
31'b0100001000100001010000000000000,
31'b0010010000000000000101000000010,
31'b1100000000000000010000100000001,
31'b1001000000000000000000010101000,
31'b0100001100000100000000000010000,
31'b0100001100000010000000000010000,
31'b0100001100000000000000000010000,
31'b1010000000000000000001100000010,
31'b1000100000100000000000000000011,
31'b0001000011000000001000001000000,
31'b0011000000001000000000101000000,
31'b0100001000010000000100000000100,
31'b1010000010100000000000010000000,
31'b0001000000000000010110000000000,
31'b0011000000000000000000101000000,
31'b0100010000000000100001000000000,
31'b0100010000000010100001000000000,
31'b0000010000000000001100010000000,
31'b1000010000000000100000000001001,
31'b0100001000000000000100000000100,
31'b0100001000000010000100000000100,
31'b0000000000000000100000001010000,
31'b0010000000100000000100000000001,
31'b1000100000000010000000000000011,
31'b1000100000000000000000000000011,
31'b0100100000000000000001000001010,
31'b0010000000000000000000000100110,
31'b1010000010000010000000010000000,
31'b1010000010000000000000010000000,
31'b0010000000000000110001000000000,
31'b0000100000000000000010000010000,
31'b0101001100000000000000000001000,
31'b1000100000010000000000000000011,
31'b1000000000000010000000010110000,
31'b1000000000000000000000010110000,
31'b0110000110000000100000000000000,
31'b0010000000000100000100000000001,
31'b0010000000000010000100000000001,
31'b0010000000000000000100000000001,
31'b1010101000000000000000000000000,
31'b0000000000000101000001000000000,
31'b0000000000000011000001000000000,
31'b0000000000000001000001000000000,
31'b1010101000001000000000000000000,
31'b0010000100010000000000001000000,
31'b0000001000010000000100000000010,
31'b0000000000001001000001000000000,
31'b1010101000010000000000000000000,
31'b0010000100001000000000001000000,
31'b0000001000001000000100000000010,
31'b0000000000010001000001000000000,
31'b0010000100000010000000001000000,
31'b0010000100000000000000001000000,
31'b0000001000000000000100000000010,
31'b0000010000000000010000000100000,
31'b0110000000000010000000000100000,
31'b0110000000000000000000000100000,
31'b0100001000000000000000100001000,
31'b0000000000100001000001000000000,
31'b0110000000001010000000000100000,
31'b0110000000001000000000000100000,
31'b0100001000001000000000100001000,
31'b0100000010010000000000000010000,
31'b0110000000010010000000000100000,
31'b0110000000010000000000000100000,
31'b0100001000010000000000100001000,
31'b0100000010001000000000000010000,
31'b0110001001000000100000000000000,
31'b0100000010000100000000000010000,
31'b0100000010000010000000000010000,
31'b0100000010000000000000000010000,
31'b1010101001000000000000000000000,
31'b0010000000000000100010010000000,
31'b0000011000000000110000000000000,
31'b0000000001000001000001000000000,
31'b0001000010000000000100100000010,
31'b0010000101010000000000001000000,
31'b0000010000000001000000000000011,
31'b0000000001001001000001000000000,
31'b1110000100000000000010000000000,
31'b0010000101001000000000001000000,
31'b0000011000010000110000000000000,
31'b0000000001010001000001000000000,
31'b0110001000100000100000000000000,
31'b0010000101000000000000001000000,
31'b0000001001000000000100000000010,
31'b0000000000000000100000000000101,
31'b0110000001000010000000000100000,
31'b0110000001000000000000000100000,
31'b0101000000000010101000000000000,
31'b0101000000000000101000000000000,
31'b1010000000000000000010001100000,
31'b1010001100000000000000010000000,
31'b1000010100000000010010000000000,
31'b0101000000001000101000000000000,
31'b0101000010000000000000000001000,
31'b0110000001010000000000000100000,
31'b1001000100000000001000010000000,
31'b1001000010000000000001000000001,
31'b0110001000000000100000000000000,
31'b0110001000000010100000000000000,
31'b0110001000000100100000000000000,
31'b0100000011000000000000000010000,
31'b1010101010000000000000000000000,
31'b0010010000000000010000000010000,
31'b0000001000000000000010010010000,
31'b0000000010000001000001000000000,
31'b1001100000000000100000000001000,
31'b0100010100000000000001000100000,
31'b0100000000110010000000000010000,
31'b0100000000110000000000000010000,
31'b0101000001100000000000000001000,
31'b0100000100000001010000000000000,
31'b0100000000101010000000000010000,
31'b0100000000101000000000000010000,
31'b0100000101000000000100000000100,
31'b0100000000100100000000000010000,
31'b0100000000100010000000000010000,
31'b0100000000100000000000000010000,
31'b0110000010000010000000000100000,
31'b0110000010000000000000000100000,
31'b0100001010000000000000100001000,
31'b0100000000011000000000000010000,
31'b0100000001000000001000100100000,
31'b0100000000010100000000000010000,
31'b0100000000010010000000000010000,
31'b0100000000010000000000000010000,
31'b0101000001000000000000000001000,
31'b0000010000000000000001001000000,
31'b0100000000001010000000000010000,
31'b0100000000001000000000000010000,
31'b0100000000000110000000000010000,
31'b0100000000000100000000000010000,
31'b0100000000000010000000000010000,
31'b0100000000000000000000000010000,
31'b0101000000110000000000000001000,
31'b1000100000000100100000000010000,
31'b1010000000000000010011000000000,
31'b1000100000000000100000000010000,
31'b0001000000000000000100100000010,
31'b1000101000000000001000100000000,
31'b0011010000000000010000000001000,
31'b1100000000000000001001000000100,
31'b0101000000100000000000000001000,
31'b0101000000100010000000000001000,
31'b1011100000000000000000100000000,
31'b1001000000100000000001000000001,
31'b0100000100000000000100000000100,
31'b0100000100000010000100000000100,
31'b0100000100000100000100000000100,
31'b0100000001100000000000000010000,
31'b0101000000010000000000000001000,
31'b0110000011000000000000000100000,
31'b1001000000000000110100000000000,
31'b1001000000010000000001000000001,
31'b0100000000000000001000100100000,
31'b0100000001010100000000000010000,
31'b0100000001010010000000000010000,
31'b0100000001010000000000000010000,
31'b0101000000000000000000000001000,
31'b0101000000000010000000000001000,
31'b1000000000000000000010001010000,
31'b1001000000000000000001000000001,
31'b0000000000000000000000001000011,
31'b0100000001000100000000000010000,
31'b0100000001000010000000000010000,
31'b0100000001000000000000000010000,
31'b1010101100000000000000000000000,
31'b0010000000011000000000001000000,
31'b0001001000000000001000001000000,
31'b0000000100000001000001000000000,
31'b0010000000010010000000001000000,
31'b0010000000010000000000001000000,
31'b0010100000000001001000000000010,
31'b0010000000010100000000001000000,
31'b1000000000000001001100000000000,
31'b0010000000001000000000001000000,
31'b1011000000000000000001000000010,
31'b0010000000001100000000001000000,
31'b0010000000000010000000001000000,
31'b0010000000000000000000001000000,
31'b0010000000000110000000001000000,
31'b0010000000000100000000001000000,
31'b0110000100000010000000000100000,
31'b0110000100000000000000000100000,
31'b0100010000000010010000001000000,
31'b0100010000000000010000001000000,
31'b0010100000000000100010000000000,
31'b0000000000000000010001000010000,
31'b1000010001000000010010000000000,
31'b0010010010000001000000000000000,
31'b1010000000000000100000010100000,
31'b0010000000101000000000001000000,
31'b1001000001000000001000010000000,
31'b0100010000010000010000001000000,
31'b0010000000100010000000001000000,
31'b0010000000100000000000001000000,
31'b0100001000000000000000001000101,
31'b0100000110000000000000000010000,
31'b1110000000010000000010000000000,
31'b0010000100000000100010010000000,
31'b0001001001000000001000001000000,
31'b0000000101000001000001000000000,
31'b0110100000000000000000010100000,
31'b0010000001010000000000001000000,
31'b1100000000000000000000010000101,
31'b0010000001010100000000001000000,
31'b1110000000000000000010000000000,
31'b0010000001001000000000001000000,
31'b1110000000000100000010000000000,
31'b0010000001001100000000001000000,
31'b0100000010000000000100000000100,
31'b0010000001000000000000001000000,
31'b0110000000000000000000000010011,
31'b0010000001000100000000001000000,
31'b0001000010000000001100000000001,
31'b1101000000000000010000000000001,
31'b0001000000000000010001000001000,
31'b0101000100000000101000000000000,
31'b1010001000000010000000010000000,
31'b1010001000000000000000010000000,
31'b1000010000000000010010000000000,
31'b1010001000000100000000010000000,
31'b1110000000100000000010000000000,
31'b0010101000000000000010000100000,
31'b1001000000000000001000010000000,
31'b1001000000000010001000010000000,
31'b0110001100000000100000000000000,
31'b0010000001100000000000001000000,
31'b1001000000001000001000010000000,
31'b0100000111000000000000000010000,
31'b0100000001000000000000000100011,
31'b0100000000010001010000000000000,
31'b0000000000000010000000001110000,
31'b0000000000000000000000001110000,
31'b0100010000000010000001000100000,
31'b0100010000000000000001000100000,
31'b1000010000000000000000000101001,
31'b0010010000100001000000000000000,
31'b0100000000000011010000000000000,
31'b0100000000000001010000000000000,
31'b0100100001000000000000010010000,
31'b0100000000000101010000000000000,
31'b0100000001000000000100000000100,
31'b0010000010000000000000001000000,
31'b0100000100100010000000000010000,
31'b0100000100100000000000000010000,
31'b1000100000000000100100000000100,
31'b0110000110000000000000000100000,
31'b1000010000000000001100001000000,
31'b0010010000001001000000000000000,
31'b1000111000000000000001000000000,
31'b0010010000000101000000000000000,
31'b1000000000000000100000010010000,
31'b0010010000000001000000000000000,
31'b0101000101000000000000000001000,
31'b0100000000100001010000000000000,
31'b0100100000000000010000000001100,
31'b0100000100001000000000000010000,
31'b0100000100000110000000000010000,
31'b0100000100000100000000000010000,
31'b0100000100000010000000000010000,
31'b0100000100000000000000000010000,
31'b0100000000000000000000000100011,
31'b0100000001010001010000000000000,
31'b0100100000010000000000010010000,
31'b0000100000000001000000100000010,
31'b0100000000010000000100000000100,
31'b0100010001000000000001000100000,
31'b1100000000000000000010000110000,
31'b0011001000000000000000101000000,
31'b0000000000000000001000101000000,
31'b0100000001000001010000000000000,
31'b0100100000000000000000010010000,
31'b0100100000000010000000010010000,
31'b0100000000000000000100000000100,
31'b0100000000000010000100000000100,
31'b0100000000000100000100000000100,
31'b0100000101100000000000000010000,
31'b0001000000000000001100000000001,
31'b1001000000000000100000010001000,
31'b0010010000000000010100000000100,
31'b0010010001001001000000000000000,
31'b0100000100000000001000100100000,
31'b1010001010000000000000010000000,
31'b1000010010000000010010000000000,
31'b0010010001000001000000000000000,
31'b0101000100000000000000000001000,
31'b0101000100000010000000000001000,
31'b1001000010000000001000010000000,
31'b1001000100000000000001000000001,
31'b0100000000100000000100000000100,
31'b0100000101000100000000000010000,
31'b0100000101000010000000000010000,
31'b0100000101000000000000000010000,
31'b1010110000000000000000000000000,
31'b1010110000000010000000000000000,
31'b0000000001000000110000000000000,
31'b0000011000000001000001000000000,
31'b1010110000001000000000000000000,
31'b0101000000000000000010000100100,
31'b0000010000010000000100000000010,
31'b0000001000010000010000000100000,
31'b1100000001000000000100000001000,
31'b0000001010100000000001001000000,
31'b0000010000001000000100000000010,
31'b0000001000001000010000000100000,
31'b0010000000000000010000100001000,
31'b0000001000000100010000000100000,
31'b0000010000000000000100000000010,
31'b0000001000000000010000000100000,
31'b1010110000100000000000000000000,
31'b1010000010000000001000000000010,
31'b0100010000000000000000100001000,
31'b0100010000000010000000100001000,
31'b1000000001000000000000100000010,
31'b1000100000000000001000010000001,
31'b1100100000010000010000000000000,
31'b0010001110000001000000000000000,
31'b0001001000000000000000010100100,
31'b0000001010000000000001001000000,
31'b1100100000001000010000000000000,
31'b0000100010001000001100000000000,
31'b1100100000000100010000000000000,
31'b0000100010000100001100000000000,
31'b1100100000000000010000000000000,
31'b0000100010000000001100000000000,
31'b0000000000000100110000000000000,
31'b1000000010000000000001010000000,
31'b0000000000000000110000000000000,
31'b0000000000000010110000000000000,
31'b1000000000100000000000100000010,
31'b1000000010001000000001010000000,
31'b0000000000001000110000000000000,
31'b0000000000001010110000000000000,
31'b1100000000000000000100000001000,
31'b0000000010000000011000000001000,
31'b0000000000010000110000000000000,
31'b0000000000000000000101000000001,
31'b1100000000001000000100000001000,
31'b0000101000000000001000001000001,
31'b0000010001000000000100000000010,
31'b0000001001000000010000000100000,
31'b1000000000001000000000100000010,
31'b1000000010100000000001010000000,
31'b0000000000100000110000000000000,
31'b0001000000000000000001101000000,
31'b1000000000000000000000100000010,
31'b1000000000000010000000100000010,
31'b1000000000000100000000100000010,
31'b1000000000000110000000100000010,
31'b1100000000100000000100000001000,
31'b0000101000000000000100000101000,
31'b0010100000000000000100100000000,
31'b0000100000000000010010001000000,
31'b1000000000010000000000100000010,
31'b1100000000000001000000010010000,
31'b1100100001000000010000000000000,
31'b0000100011000000001100000000000,
31'b1010110010000000000000000000000,
31'b1000000001000000000001010000000,
31'b0000010000000000000010010010000,
31'b1010000000000001100010000000000,
31'b1000100100100000000001000000000,
31'b1010000100000000000000100000001,
31'b0001000001000000000000011000010,
31'b0010001100100001000000000000000,
31'b0100000101000000100001000000000,
31'b0000001000100000000001001000000,
31'b0001000100000000100010000000010,
31'b0000100000101000001100000000000,
31'b0010010000000000000000000010101,
31'b0000100001000000000011000100000,
31'b0001000000000000011000000010000,
31'b0000100000100000001100000000000,
31'b1010000000000010001000000000010,
31'b1010000000000000001000000000010,
31'b0100010010000000000000100001000,
31'b1010000000000100001000000000010,
31'b1000100100000000000001000000000,
31'b1010000000001000001000000000010,
31'b1001001000010000000000000000010,
31'b0010001100000001000000000000000,
31'b0001000100000001001000000000000,
31'b0000001000000000000001001000000,
31'b1010100000000001000000001000000,
31'b0000100000001000001100000000000,
31'b1001001000000100000000000000010,
31'b0000100000000100001100000000000,
31'b1001001000000000000000000000010,
31'b0000100000000000001100000000000,
31'b1000000000000010000001010000000,
31'b1000000000000000000001010000000,
31'b0000000010000000110000000000000,
31'b1000000000000100000001010000000,
31'b1000000010100000000000100000010,
31'b1000000000001000000001010000000,
31'b0001000000000000000000011000010,
31'b1000000000001100000001010000000,
31'b0100000100000000100001000000000,
31'b0000000000000000011000000001000,
31'b0000000100000000001100010000000,
31'b0000000010000000000101000000001,
31'b0110000000000000000010000001100,
31'b0000100000000000000011000100000,
31'b0001000001000000011000000010000,
31'b0000100001100000001100000000000,
31'b1000000010001000000000100000010,
31'b1000000000100000000001010000000,
31'b0000000010100000110000000000000,
31'b1001000000000000100000000100010,
31'b1000000010000000000000100000010,
31'b1000000010000010000000100000010,
31'b1001000000000000010001000000100,
31'b0110010000000000001000000001000,
31'b0101011000000000000000000001000,
31'b0000001001000000000001001000000,
31'b0010100010000000000100100000000,
31'b0000100010000000010010001000000,
31'b1100001000000000000011000000000,
31'b0000100001000100001100000000000,
31'b1001001001000000000000000000010,
31'b0000100001000000001100000000000,
31'b1000000001000000001000000000001,
31'b1000100000000000000000110000010,
31'b0001010000000000001000001000000,
31'b0100001000100000010000001000000,
31'b1000100010100000000001000000000,
31'b1010000010000000000000100000001,
31'b0001010000001000001000001000000,
31'b0010001010100001000000000000000,
31'b1100100000000001000000000010000,
31'b0010100000000000000000100010100,
31'b0001010000010000001000001000000,
31'b1100000001000000010000010000000,
31'b0010011000000010000000001000000,
31'b0010011000000000000000001000000,
31'b0000010100000000000100000000010,
31'b0010000000000000000100110000000,
31'b1000100010001000000001000000000,
31'b0100001000000100010000001000000,
31'b0100010100000000000000100001000,
31'b0100001000000000010000001000000,
31'b1000100010000000000001000000000,
31'b1010010001000000000000010000000,
31'b1000100010000100000001000000000,
31'b0010001010000001000000000000000,
31'b0001000010000001001000000000000,
31'b0001000000000000000010001000100,
31'b0010000010000000000101000000010,
31'b1100000000000000000000000011100,
31'b1101000001000000000000000000100,
31'b0011000001000001000000100000000,
31'b1100100100000000010000000000000,
31'b0010001010010001000000000000000,
31'b1000000000000000001000000000001,
31'b1000000000000010001000000000001,
31'b0000000100000000110000000000000,
31'b0100000000000000001001000001000,
31'b1000000000001000001000000000001,
31'b1010010000100000000000010000000,
31'b0000000100001000110000000000000,
31'b0100100000000000010010000100000,
31'b1000000000010000001000000000001,
31'b1100000000000100010000010000000,
31'b0000000100010000110000000000000,
31'b1100000000000000010000010000000,
31'b1101000000100000000000000000100,
31'b0011000000100001000000100000000,
31'b0000010101000000000100000000010,
31'b1100000000001000010000010000000,
31'b1000000000100000001000000000001,
31'b1010010000001000000000010000000,
31'b0000001000000001001000100000000,
31'b0100001001000000010000001000000,
31'b0000000000000001100000000010000,
31'b1010010000000000000000010000000,
31'b1000001000000000010010000000000,
31'b1010010000000100000000010000000,
31'b1101000000001000000000000000100,
31'b0011000000001001000000100000000,
31'b0010100100000000000100100000000,
31'b1100000000100000010000010000000,
31'b1101000000000000000000000000100,
31'b0011000000000001000000100000000,
31'b1101000000000100000000000000100,
31'b0011000000000101000000100000000,
31'b1000100000101000000001000000000,
31'b1010000000001000000000100000001,
31'b0001010010000000001000001000000,
31'b0010001000101001000000000000000,
31'b1000100000100000000001000000000,
31'b1010000000000000000000100000001,
31'b1000100000100100000001000000000,
31'b0010001000100001000000000000000,
31'b0100000001000000100001000000000,
31'b0100011000000001010000000000000,
31'b0001000000000000100010000000010,
31'b1000000001000000100000000001001,
31'b1001000000000000100000000010001,
31'b1010000000010000000000100000001,
31'b0001000100000000011000000010000,
31'b0010001000110001000000000000000,
31'b1000100000001000000001000000000,
31'b1010000100000000001000000000010,
31'b1000100000001100000001000000000,
31'b0010001000001001000000000000000,
31'b1000100000000000000001000000000,
31'b1000100000000010000001000000000,
31'b1000100000000100000001000000000,
31'b0010001000000001000000000000000,
31'b0001000000000001001000000000000,
31'b0001000000000011001000000000000,
31'b0010000000000000000101000000010,
31'b0010001000011001000000000000000,
31'b1000100000010000000001000000000,
31'b1011000000000000000100001000000,
31'b1001001100000000000000000000010,
31'b0010001000010001000000000000000,
31'b1000000010000000001000000000001,
31'b1000000100000000000001010000000,
31'b0000000110000000110000000000000,
31'b1000000100000100000001010000000,
31'b1000100001100000000001000000000,
31'b1010000001000000000000100000001,
31'b0001010000000000010110000000000,
31'b0011010000000000000000101000000,
31'b0100000000000000100001000000000,
31'b0100000000000010100001000000000,
31'b0000000000000000001100010000000,
31'b1000000000000000100000000001001,
31'b0100000000001000100001000000000,
31'b0100000000001010100001000000000,
31'b0000010000000000100000001010000,
31'b1010000000000001000000011000000,
31'b1000100001001000000001000000000,
31'b1000110000000000000000000000011,
31'b0010001000000000010100000000100,
31'b0010010000000000000000000100110,
31'b1000100001000000000001000000000,
31'b1010010010000000000000010000000,
31'b1000100001000100000001000000000,
31'b0010001001000001000000000000000,
31'b0100000000100000100001000000000,
31'b0101000000000000010000101000000,
31'b0010000000000001100000000100000,
31'b1000010000000000000000010110000,
31'b1101000010000000000000000000100,
31'b0011000010000001000000100000000,
31'b0010010000000010000100000000001,
31'b0010010000000000000100000000001,
31'b1010111000000000000000000000000,
31'b0010000010000000010000000010000,
31'b0000010000000011000001000000000,
31'b0000010000000001000001000000000,
31'b0100000000000011000000001010000,
31'b0100000000000001000000001010000,
31'b0000000001000001000000000000011,
31'b0000000000010000010000000100000,
31'b0001000010000000110000100000000,
31'b0000000010100000000001001000000,
31'b0000000000001010010000000100000,
31'b0000000000001000010000000100000,
31'b0000000000000110010000000100000,
31'b0000000000000100010000000100000,
31'b0000000000000010010000000100000,
31'b0000000000000000010000000100000,
31'b0110010000000010000000000100000,
31'b0110010000000000000000000100000,
31'b0100011000000000000000100001000,
31'b0100000100000000010000001000000,
31'b1001100000000000000010000000100,
31'b0110010000001000000000000100000,
31'b1001000010010000000000000000010,
31'b0010000110000001000000000000000,
31'b0001000000000000000000010100100,
31'b0000000010000000000001001000000,
31'b1001000010001000000000000000010,
31'b0000000010000100000001001000000,
31'b1001000010000100000000000000010,
31'b0000000010001000000001001000000,
31'b1001000010000000000000000000010,
31'b0000000000100000010000000100000,
31'b1000000000000001000010000010000,
31'b1000001010000000000001010000000,
31'b0000001000000000110000000000000,
31'b0000010001000001000001000000000,
31'b0000000000000101000000000000011,
31'b0100100000000000000000100100010,
31'b0000000000000001000000000000011,
31'b0000000001010000010000000100000,
31'b1100001000000000000100000001000,
31'b0000100000100000000100000101000,
31'b0000001000010000110000000000000,
31'b0000001000000000000101000000001,
31'b0000100000000010001000001000001,
31'b0000100000000000001000001000001,
31'b0000000001000010010000000100000,
31'b0000000001000000010000000100000,
31'b1000001000001000000000100000010,
31'b0110010001000000000000000100000,
31'b0000001000100000110000000000000,
31'b0101010000000000101000000000000,
31'b1000001000000000000000100000010,
31'b1000001000000010000000100000010,
31'b1000000100000000010010000000000,
31'b1010000000000000000000000101010,
31'b0110000000000000000101000000100,
31'b0000100000000000000100000101000,
31'b0010101000000000000100100000000,
31'b0000101000000000010010001000000,
31'b1100000010000000000011000000000,
31'b0000100000100000001000001000001,
31'b1001000011000000000000000000010,
31'b0000000010000000000010000001001,
31'b0010000000000010010000000010000,
31'b0010000000000000010000000010000,
31'b0010100001000001000000010000000,
31'b0010000000000100010000000010000,
31'b0100000100000010000001000100000,
31'b0100000100000000000001000100000,
31'b1001000000110000000000000000010,
31'b0010000100100001000000000000000,
31'b0001000000000000110000100000000,
31'b0000000000100000000001001000000,
31'b1001000000101000000000000000010,
31'b0000000010001000010000000100000,
31'b1001000000100100000000000000010,
31'b0000000010000100010000000100000,
31'b1001000000100000000000000000010,
31'b0000000010000000010000000100000,
31'b0011100000000000000100000000000,
31'b0000000000010000000001001000000,
31'b1001000000011000000000000000010,
31'b0010000100001001000000000000000,
31'b1001000000010100000000000000010,
31'b0010000100000101000000000000000,
31'b1001000000010000000000000000010,
31'b0010000100000001000000000000000,
31'b0000000000000010000001001000000,
31'b0000000000000000000001001000000,
31'b1001000000001000000000000000010,
31'b0000000000000100000001001000000,
31'b1001000000000100000000000000010,
31'b0000000000001000000001001000000,
31'b1001000000000000000000000000010,
31'b0100010000000000000000000010000,
31'b1000001000000010000001010000000,
31'b1000001000000000000001010000000,
31'b0010100000000001000000010000000,
31'b1000110000000000100000000010000,
31'b0011000000000100010000000001000,
31'b1100000000000000000100100010000,
31'b0011000000000000010000000001000,
31'b0011000000000010010000000001000,
31'b0101010000100000000000000001000,
31'b0000001000000000011000000001000,
31'b0010100000010001000000010000000,
31'b0000001010000000000101000000001,
31'b1100000000100000000011000000000,
31'b0000101000000000000011000100000,
31'b1010000000000001000010000100000,
31'b0000000011000000010000000100000,
31'b0101010000010000000000000001000,
31'b0010000000000000000000010001100,
31'b0010100000100001000000010000000,
31'b0010000101001001000000000000000,
31'b1100000000010000000011000000000,
31'b0010000101000101000000000000000,
31'b1001000001010000000000000000010,
31'b0010000101000001000000000000000,
31'b0101010000000000000000000001000,
31'b0000000001000000000001001000000,
31'b1001000001001000000000000000010,
31'b0000000001000100000001001000000,
31'b1100000000000000000011000000000,
31'b0000000001001000000001001000000,
31'b1001000001000000000000000000010,
31'b0000000000000000000010000001001,
31'b1000100000000000000110000001000,
31'b0100000010001000000001000100000,
31'b0101000000000000100001100000000,
31'b0100000000100000010000001000000,
31'b0101000000000000000000011000100,
31'b0100000010000000000001000100000,
31'b1000000010000000000000000101001,
31'b0010000010100001000000000000000,
31'b1010000000000000000000000011001,
31'b0010010000001000000000001000000,
31'b0110000000000010000001000010000,
31'b0110000000000000000001000010000,
31'b0010010000000010000000001000000,
31'b0010010000000000000000001000000,
31'b0010000000000000000010000001010,
31'b0000000100000000010000000100000,
31'b0100000000000110010000001000000,
31'b0100000000000100010000001000000,
31'b0100000000000010010000001000000,
31'b0100000000000000010000001000000,
31'b1000101010000000000001000000000,
31'b0010000010000101000000000000000,
31'b1000000001000000010010000000000,
31'b0010000010000001000000000000000,
31'b0000000000000011000000000110000,
31'b0000000000000001000000000110000,
31'b0100100000000000000000100010001,
31'b0100000000010000010000001000000,
31'b0010010000100010000000001000000,
31'b0010010000100000000000001000000,
31'b1001000110000000000000000000010,
31'b0010000010010001000000000000000,
31'b1000001000000000001000000000001,
31'b1001000000000000000010010000100,
31'b0000001100000000110000000000000,
31'b0100001000000000001001000001000,
31'b1000001000001000001000000000001,
31'b0100100000000000000100001001000,
31'b1000000000100000010010000000000,
31'b1011000000010000000000000000001,
31'b1110010000000000000010000000000,
31'b0011000000000000000010000010010,
31'b0000100010000000100000100000100,
31'b1100001000000000010000010000000,
31'b0111000000000000000001000001000,
31'b0010010001000000000000001000000,
31'b1011000000000010000000000000001,
31'b1011000000000000000000000000001,
31'b0000000000000101001000100000000,
31'b0100100000000000001000000100001,
31'b0000000000000001001000100000000,
31'b0100000001000000010000001000000,
31'b1000000000000100010010000000000,
31'b1010011000000000000000010000000,
31'b1000000000000000010010000000000,
31'b1000000000000010010010000000000,
31'b0000100000000100010000010100000,
31'b0000100000000000000000101000010,
31'b0000100000000000010000010100000,
31'b0100000001010000010000001000000,
31'b1101001000000000000000000000100,
31'b0011001000000001000000100000000,
31'b1000000000010000010010000000000,
31'b1011000000100000000000000000001,
31'b0100000000001010000001000100000,
31'b0100000000001000000001000100000,
31'b1000000000100000001100001000000,
31'b0010000000101001000000000000000,
31'b0100000000000010000001000100000,
31'b0100000000000000000001000100000,
31'b1000000000000000000000000101001,
31'b0010000000100001000000000000000,
31'b0100010000000011010000000000000,
31'b0100010000000001010000000000000,
31'b1001000000000000001000100000001,
31'b0110000010000000000001000010000,
31'b0100010001000000000100000000100,
31'b0100000000010000000001000100000,
31'b1001000100100000000000000000010,
31'b0010000000110001000000000000000,
31'b1000101000001000000001000000000,
31'b0010000000001101000000000000000,
31'b1000000000000000001100001000000,
31'b0010000000001001000000000000000,
31'b1000101000000000000001000000000,
31'b0010000000000101000000000000000,
31'b0010000000000011000000000000000,
31'b0010000000000001000000000000000,
31'b0001001000000001001000000000000,
31'b0000000100000000000001001000000,
31'b1001000100001000000000000000010,
31'b0010000000011001000000000000000,
31'b1001000100000100000000000000010,
31'b0010000000010101000000000000000,
31'b1001000100000000000000000000010,
31'b0010000000010001000000000000000,
31'b1000001010000000001000000000001,
31'b1001000000000000000000000110001,
31'b0010100100000001000000010000000,
31'b0011100000000000000000000010100,
31'b0100010000010000000100000000100,
31'b0100000001000000000001000100000,
31'b1000000010100000010010000000000,
31'b0010000001100001000000000000000,
31'b0100001000000000100001000000000,
31'b0100010001000001010000000000000,
31'b0000100000000000100000100000100,
31'b1001100000000000000000010000010,
31'b0100010000000000000100000000100,
31'b0100010000000010000100000000100,
31'b0100010000000100000100000000100,
31'b1011000010000000000000000000001,
31'b0011000000000001000000000011000,
31'b0010000100000000000000010001100,
31'b0010000000000000010100000000100,
31'b0010000001001001000000000000000,
31'b1000101001000000000001000000000,
31'b0010000001000101000000000000000,
31'b1000000010000000010010000000000,
31'b0010000001000001000000000000000,
31'b0101010100000000000000000001000,
31'b0000000101000000000001001000000,
31'b0010001000000001100000000100000,
31'b0010000001011001000000000000000,
31'b1100000100000000000011000000000,
31'b0010000001010101000000000000000,
31'b1001000101000000000000000000010,
31'b0010000001010001000000000000000,
31'b1011000000000000000000000000000,
31'b1011000000000010000000000000000,
31'b1011000000000100000000000000000,
31'b1011000000000110000000000000000,
31'b1011000000001000000000000000000,
31'b1011000000001010000000000000000,
31'b1011000000001100000000000000000,
31'b1000001000010000001000000000000,
31'b1011000000010000000000000000000,
31'b0000000100000001000000000000010,
31'b1011000000010100000000000000000,
31'b1000001000001000001000000000000,
31'b1011000000011000000000000000000,
31'b1000001000000100001000000000000,
31'b1000001000000010001000000000000,
31'b1000001000000000001000000000000,
31'b1011000000100000000000000000000,
31'b1011000000100010000000000000000,
31'b1100000000000000001010010000000,
31'b0000010110000000000000001000010,
31'b1011000000101000000000000000000,
31'b0100100001000000000000100010000,
31'b0100100000010000001000000100000,
31'b0000000001000000001000011000000,
31'b1011000000110000000000000000000,
31'b1000000000000000010010000000001,
31'b0100100000001000001000000100000,
31'b0000000100000000101010000000000,
31'b0100100000000100001000000100000,
31'b0000000000000100010000000010010,
31'b0100100000000000001000000100000,
31'b0000000000000000010000000010010,
31'b1011000001000000000000000000000,
31'b1011000001000010000000000000000,
31'b1000000000000000101000000100000,
31'b1010000000001000000000000011000,
31'b1011000001001000000000000000000,
31'b1010000000000100000000000011000,
31'b1010000000000010000000000011000,
31'b1010000000000000000000000011000,
31'b1011000001010000000000000000000,
31'b1000000010000000000000000101000,
31'b1010001010000000000000100000000,
31'b1000001001001000001000000000000,
31'b0100100000000000000111000000000,
31'b1000001001000100001000000000000,
31'b1001000000000000100000100001000,
31'b1000001001000000001000000000000,
31'b1011000001100000000000000000000,
31'b0100100000001000000000100010000,
31'b1010000000000001000100010000000,
31'b0000010000000000100100000010000,
31'b0100100000000010000000100010000,
31'b0100100000000000000000100010000,
31'b0000000000000010001000011000000,
31'b0000000000000000001000011000000,
31'b0010000010000001000000000000001,
31'b1000000010100000000000000101000,
31'b0011010000000000000100100000000,
31'b0001010000000000010010001000000,
31'b0100000000000000010000001000001,
31'b0100100000010000000000100010000,
31'b0100100001000000001000000100000,
31'b0000000001000000010000000010010,
31'b1011000010000000000000000000000,
31'b1011000010000010000000000000000,
31'b1011000010000100000000000000000,
31'b0100010000000000000100000000101,
31'b1000001000000000100000000001000,
31'b1001000001000000001000100000000,
31'b1001000000010000000000000110000,
31'b1010000000000000100000100100000,
31'b1011000010010000000000000000000,
31'b1000000001000000000000000101000,
31'b1010001001000000000000100000000,
31'b1000001010001000001000000000000,
31'b1001000000000100000000000110000,
31'b1000001010000100001000000000000,
31'b1001000000000000000000000110000,
31'b1000001010000000001000000000000,
31'b0000000100000000000010000001000,
31'b0010000000000000010000000100010,
31'b0010000000000000000000111000000,
31'b0000010100000000000000001000010,
31'b0010000000000000100001000000100,
31'b0100100000000000100000000101000,
31'b0010000000001000000000111000000,
31'b0001010000010000001100000000000,
31'b0010000001000001000000000000001,
31'b1000000010000000010010000000001,
31'b0010000001000101000000000000001,
31'b0001010000001000001100000000000,
31'b0010000001001001000000000000001,
31'b0010010000000001000001000000010,
31'b1001000000100000000000000110000,
31'b0001010000000000001100000000000,
31'b1011000011000000000000000000000,
31'b1000000000010000000000000101000,
31'b1010001000010000000000100000000,
31'b1001001000000000100000000010000,
31'b1001000000000010001000100000000,
31'b1001000000000000001000100000000,
31'b0100010000000001010000000000001,
31'b1010000010000000000000000011000,
31'b1000000000000010000000000101000,
31'b1000000000000000000000000101000,
31'b1010001000000000000000100000000,
31'b1000000000000100000000000101000,
31'b1010000000000000101000000010000,
31'b1000000000001000000000000101000,
31'b1010001000001000000000100000000,
31'b1000001011000000001000000000000,
31'b0010000000010001000000000000001,
31'b1001000100000000000000000000011,
31'b0010000001000000000000111000000,
31'b0001000100001000000010000010000,
31'b0010000001000000100001000000100,
31'b1100000100000000000000001001000,
31'b0000000100000000000001001000001,
31'b0001000100000000000010000010000,
31'b0010000000000001000000000000001,
31'b1000000000100000000000000101000,
31'b0010000000000101000000000000001,
31'b1000101000000000000001000000001,
31'b0010000000001001000000000000001,
31'b1000000000101000000000000101000,
31'b0010000100000000100010100000000,
31'b0001010001000000001100000000000,
31'b0000010000000000100000000000100,
31'b0000000000010001000000000000010,
31'b0000100000000000001000001000000,
31'b0000100000000010001000001000000,
31'b0000001000000000000101000000000,
31'b0000001000000010000101000000000,
31'b0000100000001000001000001000000,
31'b1010100000000001000100000000000,
31'b0000000000000011000000000000010,
31'b0000000000000001000000000000010,
31'b0000100000010000001000001000000,
31'b0000000000000101000000000000010,
31'b0000001000010000000101000000000,
31'b0000000000001001000000000000010,
31'b1001000000000001000001001000000,
31'b1000001100000000001000000000000,
31'b0000000010000000000010000001000,
31'b0000000010000010000010000001000,
31'b0000100000100000001000001000000,
31'b0000010010000000000000001000010,
31'b0000001000100000000101000000000,
31'b0100000010000000000001000010010,
31'b0000100000101000001000001000000,
31'b0001010000000000110000010000000,
31'b0000000010010000000010000001000,
31'b0000000000100001000000000000010,
31'b0000100000000000000000000001110,
31'b0000000000000000101010000000000,
31'b0000001000110000000101000000000,
31'b0000001000000000000010100010000,
31'b0110000000000000110000000000100,
31'b0000000100000000010000000010010,
31'b0000000000000000010000000100001,
31'b0000000001010001000000000000010,
31'b0000100001000000001000001000000,
31'b0100100000000001010000100000000,
31'b0000001001000000000101000000000,
31'b0000011000010000000000000100100,
31'b0000100010000000010110000000000,
31'b1100100000000000001010000000000,
31'b0000000001000011000000000000010,
31'b0000000001000001000000000000010,
31'b0100000000000010001000010100000,
31'b0100000000000000001000010100000,
31'b0000010000000001000001000000001,
31'b0000011000000000000000000100100,
31'b0010010000000000000000100001100,
31'b1100010000000001000000000001000,
31'b0000000011000000000010000001000,
31'b1010000000000001010000000001000,
31'b0000101000000000010001000001000,
31'b0001000010001000000010000010000,
31'b0000001001100000000101000000000,
31'b1100000010000000000000001001000,
31'b0000001000000000001010000100000,
31'b0001000010000000000010000010000,
31'b0011000000000010000010000100000,
31'b0011000000000000000010000100000,
31'b1000101000000000001000010000000,
31'b0001000000000000000100010000010,
31'b1100110000000000000000000000100,
31'b0011000000001000000010000100000,
31'b1100000000000000101000001000000,
31'b0001000010010000000010000010000,
31'b0000000000100000000010000001000,
31'b0000000010010001000000000000010,
31'b0000100010000000001000001000000,
31'b0000100000000001000010000000100,
31'b0000001010000000000101000000000,
31'b0100001000010000000000010001000,
31'b0000100010001000001000001000000,
31'b0010100001000000000000101000000,
31'b0000000010000011000000000000010,
31'b0000000010000001000000000000010,
31'b0000110000000000100010000000010,
31'b0000010000000000001000000001100,
31'b0100001000000010000000010001000,
31'b0100001000000000000000010001000,
31'b1001000100000000000000000110000,
31'b1000001110000000001000000000000,
31'b0000000000000000000010000001000,
31'b0000000000000010000010000001000,
31'b0000000000000100000010000001000,
31'b0000010000000000000000001000010,
31'b0000000000001000000010000001000,
31'b0100000000000000000001000010010,
31'b0000000001000000000001001000001,
31'b0001000001000000000010000010000,
31'b0000000000010000000010000001000,
31'b0000000010100001000000000000010,
31'b0000000000010100000010000001000,
31'b0000010000010000000000001000010,
31'b0000000000011000000010000001000,
31'b0100001000100000000000010001000,
31'b0010000001000000100010100000000,
31'b0001010100000000001100000000000,
31'b0000000010000000010000000100001,
31'b1001000000100000000000000000011,
31'b0000100011000000001000001000000,
31'b0010100000001000000000101000000,
31'b0000101000000000000000001101000,
31'b1100000000100000000000001001000,
31'b0000100000000000010110000000000,
31'b0010100000000000000000101000000,
31'b1010000000000000010010000000010,
31'b1000000100000000000000000101000,
31'b1010001100000000000000100000000,
31'b1000011000000000000000010000010,
31'b0010000000000100010000000010001,
31'b1100000000000000001000000000110,
31'b0010000000000000010000000010001,
31'b0010100000010000000000101000000,
31'b0000000001000000000010000001000,
31'b1001000000000000000000000000011,
31'b0000000001000100000010000001000,
31'b0001000000001000000010000010000,
31'b0000000001001000000010000001000,
31'b1100000000000000000000001001000,
31'b0000000000000000000001001000001,
31'b0001000000000000000010000010000,
31'b0010000100000001000000000000001,
31'b1001000000010000000000000000011,
31'b0010000100000101000000000000001,
31'b0001000010000000000100010000010,
31'b0010000100001001000000000000001,
31'b1100000000010000000000001001000,
31'b0010000000000000100010100000000,
31'b0001000000010000000010000010000,
31'b1011001000000000000000000000000,
31'b1011001000000010000000000000000,
31'b1011001000000100000000000000000,
31'b1000000000011000001000000000000,
31'b0000000100000000000101000000000,
31'b1000000000010100001000000000000,
31'b1000000000010010001000000000000,
31'b1000000000010000001000000000000,
31'b1011001000010000000000000000000,
31'b1000000000001100001000000000000,
31'b1000000000001010001000000000000,
31'b1000000000001000001000000000000,
31'b1000000000000110001000000000000,
31'b1000000000000100001000000000000,
31'b1000000000000010001000000000000,
31'b1000000000000000001000000000000,
31'b0010010010000000000100000000000,
31'b0111100000000000000000000100000,
31'b0011000000000001000000100000001,
31'b1101000000000000000000000000101,
31'b1000010000000000000010000000100,
31'b1000010000000010000010000000100,
31'b1000010000000100000010000000100,
31'b1000000000110000001000000000000,
31'b0100100011000000000000000001000,
31'b1000001000000000010010000000001,
31'b1010010000000000000000010000001,
31'b1000000000101000001000000000000,
31'b1000010000010000000010000000100,
31'b1000000000100100001000000000000,
31'b1000000000100010001000000000000,
31'b1000000000100000001000000000000,
31'b1011001001000000000000000000000,
31'b0100100000000001000010000000010,
31'b1010000010010000000000100000000,
31'b1001000010000000100000000010000,
31'b1000000000000000000000100110000,
31'b1000000001010100001000000000000,
31'b1000000001010010001000000000000,
31'b1000000001010000001000000000000,
31'b1010000010000100000000100000000,
31'b1000001010000000000000000101000,
31'b1010000010000000000000100000000,
31'b1000000001001000001000000000000,
31'b1000000001000110001000000000000,
31'b1000000001000100001000000000000,
31'b1000000001000010001000000000000,
31'b1000000001000000001000000000000,
31'b0100100010010000000000000001000,
31'b0100010000000000000000001000100,
31'b0100100000000010101000000000000,
31'b0100100000000000101000000000000,
31'b1000010001000000000010000000100,
31'b0000010000000000001100100000000,
31'b0000000100000000001010000100000,
31'b0000000000000000000001000010100,
31'b0100100010000000000000000001000,
31'b0100100010000010000000000001000,
31'b1010000010100000000000100000000,
31'b1000100010000000000001000000001,
31'b0100100010001000000000000001000,
31'b1000000001100100001000000000000,
31'b1000010100000000000001100000000,
31'b1000000001100000001000000000000,
31'b1000000000001000100000000001000,
31'b1010000000000000001000000110000,
31'b1010000001010000000000100000000,
31'b1001000001000000100000000010000,
31'b1000000000000000100000000001000,
31'b1000000000000010100000000001000,
31'b1000000000000100100000000001000,
31'b1000000010010000001000000000000,
31'b1010000001000100000000100000000,
31'b1000001001000000000000000101000,
31'b1010000001000000000000100000000,
31'b1000000010001000001000000000000,
31'b1000000000010000100000000001000,
31'b1000000010000100001000000000000,
31'b0100000000000000010100000000000,
31'b1000000010000000001000000000000,
31'b0010010000000000000100000000000,
31'b0010010000000010000100000000000,
31'b0010010000000100000100000000000,
31'b0010010000000110000100000000000,
31'b1000000000100000100000000001000,
31'b1000010000000001001000001000000,
31'b1000110000010000000000000000010,
31'b1000100000000001100000000000100,
31'b0100100001000000000000000001000,
31'b0101000000000000000100010000100,
31'b1010000001100000000000100000000,
31'b1000100001000000000001000000001,
31'b1000110000000100000000000000010,
31'b1000100000000000000010001001000,
31'b1000110000000000000000000000010,
31'b1000000010100000001000000000000,
31'b1010000000010100000000100000000,
31'b1001000000000100100000000010000,
31'b1010000000010000000000100000000,
31'b1001000000000000100000000010000,
31'b1000000001000000100000000001000,
31'b1001001000000000001000100000000,
31'b1010000000011000000000100000000,
31'b1001000000001000100000000010000,
31'b1010000000000100000000100000000,
31'b1000001000000000000000000101000,
31'b1010000000000000000000100000000,
31'b0100000000000001000000000000100,
31'b1010000000001100000000100000000,
31'b1000001000001000000000000101000,
31'b1010000000001000000000100000000,
31'b1000000011000000001000000000000,
31'b0100100000010000000000000001000,
31'b0100100000010010000000000001000,
31'b1010000000110000000000100000000,
31'b1001000000100000100000000010000,
31'b1100010000000000010000100000000,
31'b0010010000000001010000000000100,
31'b0001000000000011001000000000001,
31'b0001000000000001001000000000001,
31'b0100100000000000000000000001000,
31'b0100100000000010000000000001000,
31'b1010000000100000000000100000000,
31'b1000100000000000000001000000001,
31'b0100100000001000000000000001000,
31'b0100100000001010000000000001000,
31'b1010000000101000000000100000000,
31'b1000100000001000000001000000001,
31'b0000000000001000000101000000000,
31'b0000001000010001000000000000010,
31'b0000101000000000001000001000000,
31'b1001000000000000000100001000010,
31'b0000000000000000000101000000000,
31'b0000000000000010000101000000000,
31'b0000000000000100000101000000000,
31'b1000000100010000001000000000000,
31'b0000001000000011000000000000010,
31'b0000001000000001000000000000010,
31'b1010100000000000000001000000010,
31'b1000000100001000001000000000000,
31'b0000000000010000000101000000000,
31'b0000000000000000110000000000001,
31'b1000000100000010001000000000000,
31'b1000000100000000001000000000000,
31'b0000001010000000000010000001000,
31'b0000001010000010000010000001000,
31'b0000101000100000001000001000000,
31'b1100000000000000001000001100000,
31'b0000000000100000000101000000000,
31'b0000000000100010000101000000000,
31'b0000000001000000001010000100000,
31'b1000000100110000001000000000000,
31'b0100000010000001000100000010000,
31'b0000001000100001000000000000010,
31'b1000100001000000001000010000000,
31'b1000000000000000000000100000011,
31'b0000000000110000000101000000000,
31'b0000000000000000000010100010000,
31'b1000010001000000000001100000000,
31'b1000000100100000001000000000000,
31'b0000001000000000010000000100001,
31'b0000010000000000000100000000011,
31'b0000101001000000001000001000000,
31'b0010010010000000000000000010100,
31'b0000000001000000000101000000000,
31'b0000010000010000000000000100100,
31'b0000000001000100000101000000000,
31'b1000010000000000000110000010000,
31'b0000010000001010000000000100100,
31'b0000010000001000000000000100100,
31'b1010000110000000000000100000000,
31'b1000010010000000000000010000010,
31'b0000010000000010000000000100100,
31'b0000010000000000000000000100100,
31'b1000010000100000000001100000000,
31'b1000000101000000001000000000000,
31'b0000100010000000001100000000001,
31'b1100100000000000010000000000001,
31'b0000100000000000010001000001000,
31'b0110000000000000010000000100100,
31'b0000000001100000000101000000000,
31'b0000010100000000001100100000000,
31'b0000000000000000001010000100000,
31'b0000000100000000000001000010100,
31'b1100000000000000000000101010000,
31'b0011001000000000000010000100000,
31'b1000100000000000001000010000000,
31'b1000100000000010001000010000000,
31'b1000010000000100000001100000000,
31'b0000010000100000000000000100100,
31'b1000010000000000000001100000000,
31'b1000010000000010000001100000000,
31'b0000001000100000000010000001000,
31'b0100000000011000000000010001000,
31'b0000101010000000001000001000000,
31'b0010010001000000000000000010100,
31'b0000000010000000000101000000000,
31'b0100000000010000000000010001000,
31'b0000000010000100000101000000000,
31'b1000000110010000001000000000000,
31'b0100000000100001000100000010000,
31'b0100000000001000000000010001000,
31'b1010000101000000000000100000000,
31'b1000010001000000000000010000010,
31'b0100000000000010000000010001000,
31'b0100000000000000000000010001000,
31'b1000000000000000000001010000001,
31'b1000000110000000001000000000000,
31'b0000001000000000000010000001000,
31'b0000001000000010000010000001000,
31'b0000001000000100000010000001000,
31'b0010000000000000000010100100000,
31'b0000001000001000000010000001000,
31'b0100001000000000000001000010010,
31'b0000001001000000000001001000001,
31'b0011110000000001000000000000000,
31'b0100000000000001000100000010000,
31'b0100000000101000000000010001000,
31'b0101000000000000010000000001100,
31'b1010010000000000001001000000000,
31'b0100000000100010000000010001000,
31'b0100000000100000000000010001000,
31'b1000110100000000000000000000010,
31'b1010100000000000000000110000000,
31'b0000100000100000001100000000001,
31'b0010010000000100000000000010100,
31'b1010000100010000000000100000000,
31'b0010010000000000000000000010100,
31'b0000100000000000000000001101000,
31'b0110000000000000000001001000100,
31'b0000101000000000010110000000000,
31'b0010101000000000000000101000000,
31'b1010000100000100000000100000000,
31'b1000010000000100000000010000010,
31'b1010000100000000000000100000000,
31'b1000010000000000000000010000010,
31'b0101100000000000000100000000100,
31'b0100000001000000000000010001000,
31'b1010000100001000000000100000000,
31'b1000010000001000000000010000010,
31'b0000100000000000001100000000001,
31'b1001001000000000000000000000011,
31'b0000100010000000010001000001000,
31'b0010010000100000000000000010100,
31'b0000100000100000000000001101000,
31'b1100001000000000000000001001000,
31'b0000001000000000000001001000001,
31'b0001001000000000000010000010000,
31'b0100100100000000000000000001000,
31'b0100100100000010000000000001000,
31'b1010000100100000000000100000000,
31'b1000100100000000000001000000001,
31'b0100100100001000000000000001000,
31'b0100000000000000010000000010100,
31'b1010000000000000001000000000011,
31'b0101000000000001000100000001000,
31'b0000000100000000100000000000100,
31'b0110000000000000000000000010010,
31'b0010000001000000000000001000001,
31'b0110000000000100000000000010010,
31'b0010000000000000000011000001000,
31'b0110000000001000000000000010010,
31'b0010000001001000000000001000001,
31'b1110000000000000000010000000001,
31'b0010000000000001000000110000000,
31'b1100000000000000000000010000100,
31'b0010000001010000000000001000001,
31'b1100000000000100000000010000100,
31'b0010000000010000000011000001000,
31'b1100000000001000000000010000100,
31'b1101000000100000010000000000000,
31'b1000011000000000001000000000000,
31'b0010001010000000000100000000000,
31'b0110000000100000000000000010010,
31'b0010001010000100000100000000000,
31'b0000000110000000000000001000010,
31'b1000001000000000000010000000100,
31'b1001000000000000001000010000001,
31'b1101000000010000010000000000000,
31'b0001000100000000110000010000000,
31'b0010001010010000000100000000000,
31'b1100000000100000000000010000100,
31'b1101000000001000010000000000000,
31'b0001000010001000001100000000000,
31'b1101000000000100010000000000000,
31'b0010000010000001000001000000010,
31'b1101000000000000010000000000000,
31'b0001000010000000001100000000000,
31'b0010000000000100000000001000001,
31'b0110000001000000000000000010010,
31'b0010000000000000000000001000001,
31'b0010000000000010000000001000001,
31'b0010000001000000000011000001000,
31'b0000100010000000010000100100000,
31'b0010000000001000000000001000001,
31'b1010010000000000000000000011000,
31'b0010000001000001000000110000000,
31'b1100000001000000000000010000100,
31'b0010000000010000000000001000001,
31'b0010100000000000010000100010000,
31'b0000000100000001000001000000001,
31'b0000001100000000000000000100100,
31'b0010000100000000000000100001100,
31'b1100000100000001000000000001000,
31'b0100001000000010000000001000100,
31'b0100001000000000000000001000100,
31'b0010000000100000000000001000001,
31'b0000000000000000100100000010000,
31'b1001100000000000000000100000010,
31'b0000100000000000100000010000100,
31'b0010000000101000000000001000001,
31'b0000010000000000001000011000000,
31'b0011000000000100000100100000000,
31'b1100000000000000010000000011000,
31'b0011000000000000000100100000000,
31'b0001000000000000010010001000000,
31'b1100100100000000000000000000100,
31'b0010100100000001000000100000000,
31'b1101000001000000010000000000000,
31'b0001000011000000001100000000000,
31'b0010001000100000000100000000000,
31'b0110000010000000000000000010010,
31'b0100001001000000100000000000010,
31'b0100000000000000000100000000101,
31'b1001000100100000000001000000000,
31'b0100100000000000000000010010001,
31'b0100000001000001010000000000001,
31'b0100000000010000000000000100010,
31'b0010001000110000000100000000000,
31'b1100000010000000000000010000100,
31'b0100000000001010000000000100010,
31'b0100000000001000000000000100010,
31'b0100000000000110000000000100010,
31'b0100000000000100000000000100010,
31'b0100000000000010000000000100010,
31'b0100000000000000000000000100010,
31'b0010001000000000000100000000000,
31'b0010001000000010000100000000000,
31'b0010001000000100000100000000000,
31'b0000000100000000000000001000010,
31'b1001000100000000000001000000000,
31'b1001000100000010000001000000000,
31'b1001000100000100000001000000000,
31'b0001000000010000001100000000000,
31'b0010001000010000000100000000000,
31'b0010001000010010000100000000000,
31'b1011000000000001000000001000000,
31'b0001000000001000001100000000000,
31'b1001000100010000000001000000000,
31'b0010000000000001000001000000010,
31'b1000101000000000000000000000010,
31'b0001000000000000001100000000000,
31'b0100001000000100100000000000010,
31'b1001100000000000000001010000000,
31'b0100001000000000100000000000010,
31'b0100001000000010100000000000010,
31'b0100000000000101010000000000001,
31'b0000100000000000010000100100000,
31'b0100000000000001010000000000001,
31'b0100000001010000000000000100010,
31'b1010000000000000000100011000000,
31'b1000010000000000000000000101000,
31'b1010011000000000000000100000000,
31'b1000010000000100000000000101000,
31'b0000000000000011001000010000000,
31'b0000000000000001001000010000000,
31'b0100000001000010000000000100010,
31'b0100000001000000000000000100010,
31'b0100000100000000000000000010001,
31'b0100001010000000000000001000100,
31'b0100001000100000100000000000010,
31'b0000000101000000000000001000010,
31'b1100001000000000010000100000000,
31'b0010001000000001010000000000100,
31'b1100000100000000000010000000010,
31'b0001010100000000000010000010000,
31'b0010010000000001000000000000001,
31'b1000010000100000000000000101000,
31'b0011000010000000000100100000000,
31'b0001000010000000010010001000000,
31'b0010010000001001000000000000001,
31'b0010000000000000100100000100000,
31'b1001000000000000000010100000100,
31'b0001000001000000001100000000000,
31'b0000000000000000100000000000100,
31'b0000000000000010100000000000100,
31'b0000000000000100100000000000100,
31'b0000000010100000000000001000010,
31'b0000000000001000100000000000100,
31'b0000000000001010100000000000100,
31'b0000000000001100100000000000100,
31'b0001000010000000000000100100100,
31'b0000000000010000100000000000100,
31'b0000010000000001000000000000010,
31'b0000000000010100100000000000100,
31'b0000010000000101000000000000010,
31'b0000000001000001000001000000001,
31'b0000010000001001000000000000010,
31'b0010000001000000000000100001100,
31'b1100000001000001000000000001000,
31'b0000000000100000100000000000100,
31'b0000000010000100000000001000010,
31'b0000000010000010000000001000010,
31'b0000000010000000000000001000010,
31'b1001000010000000000001000000000,
31'b1001000010000010000001000000000,
31'b1001000010000100000001000000000,
31'b0001000000000000110000010000000,
31'b0000100010000001001000000000000,
31'b0000100000000000000010001000100,
31'b0000110000000000000000000001110,
31'b0000010000000000101010000000000,
31'b1100100001000000000000000000100,
31'b0010100001000001000000100000000,
31'b1101000100000000010000000000000,
31'b0001000110000000001100000000000,
31'b0000000001000000100000000000100,
31'b0000001000000000000100000000011,
31'b0010000100000000000000001000001,
31'b0010001010000000000000000010100,
31'b0000000001001000100000000000100,
31'b0000001000010000000000000100100,
31'b0010000100001000000000001000001,
31'b1100000000010001000000000001000,
31'b0000000001010000100000000000100,
31'b0000010001000001000000000000010,
31'b0010000100010000000000001000001,
31'b1100000000001001000000000001000,
31'b0000000000000001000001000000001,
31'b0000001000000000000000000100100,
31'b0010000000000000000000100001100,
31'b1100000000000001000000000001000,
31'b0100000010000000000000000010001,
31'b0100001100000000000000001000100,
31'b0110000000000000000100000000110,
31'b0000000100000000100100000010000,
31'b1100100000010000000000000000100,
31'b0010100000010001000000100000000,
31'b1100000010000000000010000000010,
31'b0001010010000000000010000010000,
31'b1100100000001000000000000000100,
31'b0011010000000000000010000100000,
31'b1100000000000000000100010010000,
31'b0001010000000000000100010000010,
31'b1100100000000000000000000000100,
31'b0010100000000001000000100000000,
31'b1000001000000000000001100000000,
31'b1100000000100001000000000001000,
31'b0000000010000000100000000000100,
31'b0000000010000010100000000000100,
31'b0000000010000100100000000000100,
31'b0000000000100000000000001000010,
31'b1001000000100000000001000000000,
31'b1001000000100010000001000000000,
31'b1001000000100100000001000000000,
31'b0001000000000000000000100100100,
31'b0000100000100001001000000000000,
31'b0000010010000001000000000000010,
31'b0000100000000000100010000000010,
31'b0000000000000000001000000001100,
31'b1001000000110000000001000000000,
31'b0100011000000000000000010001000,
31'b0110000000000000010010000001000,
31'b0100000100000000000000000100010,
31'b0000010000000000000010000001000,
31'b0000000000000100000000001000010,
31'b0000000000000010000000001000010,
31'b0000000000000000000000001000010,
31'b1001000000000000000001000000000,
31'b1001000000000010000001000000000,
31'b1001000000000100000001000000000,
31'b0000000000001000000000001000010,
31'b0000100000000001001000000000000,
31'b0000100000000011001000000000000,
31'b0000100000000101001000000000000,
31'b0000000000010000000000001000010,
31'b1001000000010000000001000000000,
31'b1010100000000000000100001000000,
31'b1001000000010100000001000000000,
31'b0001000100000000001100000000000,
31'b0100000000100000000000000010001,
31'b0110000000000000100100001000000,
31'b0100001100000000100000000000010,
31'b0010001000000000000000000010100,
31'b1100000000000001101000000000000,
31'b0010101000000000000100010000000,
31'b1100000000100000000010000000010,
31'b0010110000000000000000101000000,
31'b0101100000000000100001000000000,
31'b1000010100000000000000000101000,
31'b1000001000000010000000010000010,
31'b1000001000000000000000010000010,
31'b0001000000000000001000000010100,
31'b0000001010000000000000000100100,
31'b0010010000000000010000000010001,
31'b1100000010000001000000000001000,
31'b0100000000000000000000000010001,
31'b0100000000000010000000000010001,
31'b0100000000000100000000000010001,
31'b0000000001000000000000001000010,
31'b1001000001000000000001000000000,
31'b1100010000000000000000001001000,
31'b1100000000000000000010000000010,
31'b0001010000000000000010000010000,
31'b0100000000010000000000000010001,
31'b0100100000000000010000101000000,
31'b0100100000000000000000010100010,
31'b0000000001010000000000001000010,
31'b1100100010000000000000000000100,
31'b0010100010000001000000100000000,
31'b1100000000010000000010000000010,
31'b0001010000010000000010000010000,
31'b0010000010100000000100000000000,
31'b0110001000000000000000000010010,
31'b0100000100000000000100001010000,
31'b1001000000000000010010010000000,
31'b1000000000100000000010000000100,
31'b1000010000010100001000000000000,
31'b1000010000010010001000000000000,
31'b1000010000010000001000000000000,
31'b0010001000000001000000110000000,
31'b1100001000000000000000010000100,
31'b1010000000100000000000010000001,
31'b1000010000001000001000000000000,
31'b1000010000000110001000000000000,
31'b1000010000000100001000000000000,
31'b1000010000000010001000000000000,
31'b1000010000000000001000000000000,
31'b0010000010000000000100000000000,
31'b0100000001000000000000001000100,
31'b0010000010000100000100000000000,
31'b0110000100000000100000000000001,
31'b1000000000000000000010000000100,
31'b1000000000000010000010000000100,
31'b1000000000000100000010000000100,
31'b1000010000110000001000000000000,
31'b0010000010010000000100000000000,
31'b0110000000000000000001010001000,
31'b1010000000000000000000010000001,
31'b1010000000000010000000010000001,
31'b1000000000010000000010000000100,
31'b1000010000100100001000000000000,
31'b0000000000000000000100000110000,
31'b1000010000100000001000000000000,
31'b0100000010000100100000000000010,
31'b0100000000100000000000001000100,
31'b0100000010000000100000000000010,
31'b0100000010000010100000000000010,
31'b1000010000000000000000100110000,
31'b0000000100010000000000000100100,
31'b0101000000000000010000011000000,
31'b1000010001010000001000000000000,
31'b0100100000000000100010000000100,
31'b0100000000000000001000000001010,
31'b1010010010000000000000100000000,
31'b1000010001001000001000000000000,
31'b0000000100000010000000000100100,
31'b0000000100000000000000000100100,
31'b1000010001000010001000000000000,
31'b1000010001000000001000000000000,
31'b0100000000000010000000001000100,
31'b0100000000000000000000001000100,
31'b0100000010100000100000000000010,
31'b0100000000000100000000001000100,
31'b1000000001000000000010000000100,
31'b0000000000000000001100100000000,
31'b1000000100010000000001100000000,
31'b0000010000000000000001000010100,
31'b0100110010000000000000000001000,
31'b0100000000010000000000001000100,
31'b1010000001000000000000010000001,
31'b0100000000010100000000001000100,
31'b1000000100000100000001100000000,
31'b0000000100100000000000000100100,
31'b1000000100000000000001100000000,
31'b1000010001100000001000000000000,
31'b0010000000100000000100000000000,
31'b0010000000100010000100000000000,
31'b0100000001000000100000000000010,
31'b0100001000000000000100000000101,
31'b1000010000000000100000000001000,
31'b1000010000000010100000000001000,
31'b1000100000110000000000000000010,
31'b1000010010010000001000000000000,
31'b0010000000110000000100000000000,
31'b0010000000110010000100000000000,
31'b1010010001000000000000100000000,
31'b1000010010001000001000000000000,
31'b1000100000100100000000000000010,
31'b1000010010000100001000000000000,
31'b1000100000100000000000000000010,
31'b1000010010000000001000000000000,
31'b0010000000000000000100000000000,
31'b0010000000000010000100000000000,
31'b0010000000000100000100000000000,
31'b0010000000000110000100000000000,
31'b0010000000001000000100000000000,
31'b1000000000000001001000001000000,
31'b1000100000010000000000000000010,
31'b1000100000010010000000000000010,
31'b0010000000010000000100000000000,
31'b0010000000010010000100000000000,
31'b1000100000001000000000000000010,
31'b1010000100000000001001000000000,
31'b1000100000000100000000000000010,
31'b1000100000000110000000000000010,
31'b1000100000000000000000000000010,
31'b1000100000000010000000000000010,
31'b0100000000000100100000000000010,
31'b0100000010100000000000001000100,
31'b0100000000000000100000000000010,
31'b0100000000000010100000000000010,
31'b1100000000100000010000100000000,
31'b0010100100000000000100010000000,
31'b0100000000001000100000000000010,
31'b0100000000001010100000000000010,
31'b1010010000000100000000100000000,
31'b1000011000000000000000000101000,
31'b1010010000000000000000100000000,
31'b1000000100000000000000010000010,
31'b0001000100000000000001011000000,
31'b0000001000000001001000010000000,
31'b1010010000001000000000100000000,
31'b1000010011000000001000000000000,
31'b0010000001000000000100000000000,
31'b0100000010000000000000001000100,
31'b0100000000100000100000000000010,
31'b0100000010000100000000001000100,
31'b1100000000000000010000100000000,
31'b0010000000000001010000000000100,
31'b1100000000000100010000100000000,
31'b0011000000000000000100000011000,
31'b0100110000000000000000000001000,
31'b0100110000000010000000000001000,
31'b1010010000100000000000100000000,
31'b1000110000000000000001000000001,
31'b1100000000010000010000100000000,
31'b0010001000000000100100000100000,
31'b1000100001000000000000000000010,
31'b1000100001000010000000000000010,
31'b0000001000000000100000000000100,
31'b0000001000000010100000000000100,
31'b0100000000000000000100001010000,
31'b0110000000100000100000000000001,
31'b0000010000000000000101000000000,
31'b0000010000000010000101000000000,
31'b0000010000000100000101000000000,
31'b1000010100010000001000000000000,
31'b0000001000010000100000000000100,
31'b0000011000000001000000000000010,
31'b0101000000000000110010000000000,
31'b1000010100001000001000000000000,
31'b0000010000010000000101000000000,
31'b0000000001000000000000000100100,
31'b1000010100000010001000000000000,
31'b1000010100000000001000000000000,
31'b0010000110000000000100000000000,
31'b0110000000000100100000000000001,
31'b0110000000000010100000000000001,
31'b0110000000000000100000000000001,
31'b1000000100000000000010000000100,
31'b1000000100000010000010000000100,
31'b1000000100000100000010000000100,
31'b0110000000001000100000000000001,
31'b0010000110010000000100000000000,
31'b0001100000000001000000000110000,
31'b1010000100000000000000010000001,
31'b1010000010000000001001000000000,
31'b1000000100010000000010000000100,
31'b0000010000000000000010100010000,
31'b1000000001000000000001100000000,
31'b1000010100100000001000000000000,
31'b0000001001000000100000000000100,
31'b0000000000000000000100000000011,
31'b0100000110000000100000000000010,
31'b0010000010000000000000000010100,
31'b0000010001000000000101000000000,
31'b0000000000010000000000000100100,
31'b1000000000110000000001100000000,
31'b1000000000000000000110000010000,
31'b0000000000001010000000000100100,
31'b0000000000001000000000000100100,
31'b1000000010000010000000010000010,
31'b1000000010000000000000010000010,
31'b0000000000000010000000000100100,
31'b0000000000000000000000000100100,
31'b1000000000100000000001100000000,
31'b0000000000000100000000000100100,
31'b0100001010000000000000000010001,
31'b0100000100000000000000001000100,
31'b1000000000011000000001100000000,
31'b0110000001000000100000000000001,
31'b1000000101000000000010000000100,
31'b0000000100000000001100100000000,
31'b1000000000010000000001100000000,
31'b1000000000100000000110000010000,
31'b1000000000001100000001100000000,
31'b0001000000000000000000101000010,
31'b1000000000001000000001100000000,
31'b1000000010100000000000010000010,
31'b1000000000000100000001100000000,
31'b0000000000100000000000000100100,
31'b1000000000000000000001100000000,
31'b1000000000000010000001100000000,
31'b0010000100100000000100000000000,
31'b0010000100100010000100000000000,
31'b0100000101000000100000000000010,
31'b0010000001000000000000000010100,
31'b0011000000000000000000000001100,
31'b0101100000000000000001000100000,
31'b0011000000000100000000000001100,
31'b0011100000100001000000000000000,
31'b0010000100110000000100000000000,
31'b1100000000000001001000000100000,
31'b1000100000000000001000100000001,
31'b1000000001000000000000010000010,
31'b0110000000000000000100001100000,
31'b0100010000000000000000010001000,
31'b1000100100100000000000000000010,
31'b1000010110000000001000000000000,
31'b0010000100000000000100000000000,
31'b0010000100000010000100000000000,
31'b0010000100000100000100000000000,
31'b0000001000000000000000001000010,
31'b1001001000000000000001000000000,
31'b1001001000000010000001000000000,
31'b1001001000000100000001000000000,
31'b0011100000000001000000000000000,
31'b0010000100010000000100000000000,
31'b1010000000000100001001000000000,
31'b1010000000000010001001000000000,
31'b1010000000000000001001000000000,
31'b1001001000010000000001000000000,
31'b0100010000100000000000010001000,
31'b1000100100000000000000000000010,
31'b1010000000001000001001000000000,
31'b0100001000100000000000000010001,
31'b0010000000000100000000000010100,
31'b0100000100000000100000000000010,
31'b0010000000000000000000000010100,
31'b0011000001000000000000000001100,
31'b0010100000000000000100010000000,
31'b0100000100001000100000000000010,
31'b0010000000001000000000000010100,
31'b1000000000000110000000010000010,
31'b1000000000000100000000010000010,
31'b1000000000000010000000010000010,
31'b1000000000000000000000010000010,
31'b0001000000000000000001011000000,
31'b0000000010000000000000000100100,
31'b1000000010100000000001100000000,
31'b1000000000001000000000010000010,
31'b0100001000000000000000000010001,
31'b0100001000000010000000000010001,
31'b0100001000000100000000000010001,
31'b0010000000100000000000000010100,
31'b1100000100000000010000100000000,
31'b0010100000100000000100010000000,
31'b1100001000000000000010000000010,
31'b0011100001000001000000000000000,
31'b0100110100000000000000000001000,
31'b1001000000000000100001000100000,
31'b1000000010001000000001100000000,
31'b1000000000100000000000010000010,
31'b1001000000000000010000000000110,
31'b0000000010100000000000000100100,
31'b1000000010000000000001100000000,
31'b1000000010000010000001100000000,
31'b1011100000000000000000000000000,
31'b1011100000000010000000000000000,
31'b0000000100000000001000001000000,
31'b0001001000000001000001000000000,
31'b1011100000001000000000000000000,
31'b0100010000000000000010000100100,
31'b0001000000010000000100000000010,
31'b1010000100000001000100000000000,
31'b1011100000010000000000000000000,
31'b1000000000000000000101001000000,
31'b0001000000001000000100000000010,
31'b1000101000001000001000000000000,
31'b0010000000000001001001000000000,
31'b1000101000000100001000000000000,
31'b0001000000000000000100000000010,
31'b1000101000000000001000000000000,
31'b1011100000100000000000000000000,
31'b1010000000000000010100000010000,
31'b0101000000000000000000100001000,
31'b0101000000000010000000100001000,
31'b0100000001000010000000100010000,
31'b0100000001000000000000100010000,
31'b0100000000010000001000000100000,
31'b0100000001000100000000100010000,
31'b0100001011000000000000000001000,
31'b1000100000000000010010000000001,
31'b0100000000001000001000000100000,
31'b0110000000000000100000000011000,
31'b0100000000000100001000000100000,
31'b0100000001010000000000100010000,
31'b0100000000000000001000000100000,
31'b0100000000000010001000000100000,
31'b1011100001000000000000000000000,
31'b0100001000000001000010000000010,
31'b0001010000000000110000000000000,
31'b0100001000100000101000000000000,
31'b0100000000100010000000100010000,
31'b0100000000100000000000100010000,
31'b0001010000001000110000000000000,
31'b1100000100000000001010000000000,
31'b0100001010100000000000000001000,
31'b0000000010000001000001100000000,
31'b0001010000010000110000000000000,
31'b0010010000000000010000100010000,
31'b0100000000000000000111000000000,
31'b0100000000110000000000100010000,
31'b0001000001000000000100000000010,
31'b1000101001000000001000000000000,
31'b0100001010010000000000000001000,
31'b0100000000001000000000100010000,
31'b0101000001000000000000100001000,
31'b0100001000000000101000000000000,
31'b0100000000000010000000100010000,
31'b0100000000000000000000100010000,
31'b0100000001010000001000000100000,
31'b0100000000000100000000100010000,
31'b0100001010000000000000000001000,
31'b0100001010000010000000000001000,
31'b1000001100000000001000010000000,
31'b1000001010000000000001000000001,
31'b0000000000000001000000010000010,
31'b0100000000010000000000100010000,
31'b0100000001000000001000000100000,
31'b0100000001000010001000000100000,
31'b1100000000000000000000011001000,
31'b0000000100010000100000001001000,
31'b0001000000000000000010010010000,
31'b0000000100000001000010000000100,
31'b1001000000000000000000010000011,
31'b0000000001000000000010010001000,
31'b0001000010010000000100000000010,
31'b0010000101000000000000101000000,
31'b0100001001100000000000000001000,
31'b0000000100000000100000001001000,
31'b0001000010001000000100000000010,
31'b0010000001000000000000000001101,
31'b0011000000000000000000000010101,
31'b0010000100000001000000010000001,
31'b0001000010000000000100000000010,
31'b1000101010000000001000000000000,
31'b0110000000000000001000000010000,
31'b0110000000000010001000000010000,
31'b0110000000000100001000000010000,
31'b1000010000000001000101000000000,
31'b0110000000001000001000000010000,
31'b0100000000000000100000000101000,
31'b1000011000010000000000000000010,
31'b1000001000000001100000000000100,
31'b0100001001000000000000000001000,
31'b0101000000000000101000100000000,
31'b1000011000001000000000000000010,
31'b1000001001000000000001000000001,
31'b1000011000000100000000000000010,
31'b1000001000000000000010001001000,
31'b1000011000000000000000000000010,
31'b1000000000000000010100000100000,
31'b0100001000110000000000000001000,
31'b0000000000010001000001100000000,
31'b0001010010000000110000000000000,
31'b0010000100001000000000101000000,
31'b0000001000000000000100100000010,
31'b0000000000000000000010010001000,
31'b0000010000000000000000011000010,
31'b0010000100000000000000101000000,
31'b0100001000100000000000000001000,
31'b0000000000000001000001100000000,
31'b1010101000000000000000100000000,
31'b0010000000000000000000000001101,
31'b0100001000101000000000000001000,
31'b0000000000010000000010010001000,
31'b0001000100000000100000001010000,
31'b0010000100010000000000101000000,
31'b0100001000010000000000000001000,
31'b0100001000010010000000000001000,
31'b1000001000000000110100000000000,
31'b1000010000000000100000000100010,
31'b0100001000011000000000000001000,
31'b0100000010000000000000100010000,
31'b1000010000000000010001000000100,
31'b0111000000000000001000000001000,
31'b0100001000000000000000000001000,
31'b0100001000000010000000000001000,
31'b1000000000000001000000000100100,
31'b1000001000000000000001000000001,
31'b0100001000001000000000000001000,
31'b0100001000001010000000000001000,
31'b1000011001000000000000000000010,
31'b1000001000001000000001000000001,
31'b0000000000000100001000001000000,
31'b0000100000010001000000000000010,
31'b0000000000000000001000001000000,
31'b0000000000000010001000001000000,
31'b0000101000000000000101000000000,
31'b1010000000000101000100000000000,
31'b0000000000001000001000001000000,
31'b1010000000000001000100000000000,
31'b0000100000000011000000000000010,
31'b0000100000000001000000000000010,
31'b0000000000010000001000001000000,
31'b0000100000000101000000000000010,
31'b0011001000000010000000001000000,
31'b0011001000000000000000001000000,
31'b0001000100000000000100000000010,
31'b1010000000010001000100000000000,
31'b0000100010000000000010000001000,
31'b0000100010000010000010000001000,
31'b0000000000100000001000001000000,
31'b0000010000000001100000000001000,
31'b0000101000100000000101000000000,
31'b1100000000000000000101000100000,
31'b0000000000101000001000001000000,
31'b1010000000100001000100000000000,
31'b0000010010000001001000000000000,
31'b0000100000100001000000000000010,
31'b0000000000000000000000000001110,
31'b0000100000000000101010000000000,
31'b1100010001000000000000000000100,
31'b0011001000100000000000001000000,
31'b0100000100000000001000000100000,
31'b0100000100000010001000000100000,
31'b0000100000000000010000000100001,
31'b0100000000000101010000100000000,
31'b0000000001000000001000001000000,
31'b0100000000000001010000100000000,
31'b0000101001000000000101000000000,
31'b1100000000000100001010000000000,
31'b0000000010000000010110000000000,
31'b1100000000000000001010000000000,
31'b0000100001000011000000000000010,
31'b0000100001000001000000000000010,
31'b0000000001010000001000001000000,
31'b0100100000000000001000010100000,
31'b1100010000100000000000000000100,
31'b0011001001000000000000001000000,
31'b0001000101000000000100000000010,
31'b1100000000010000001010000000000,
31'b0000100011000000000010000001000,
31'b1100001000000000010000000000001,
31'b0000001000000000010001000001000,
31'b0100001100000000101000000000000,
31'b1100010000010000000000000000100,
31'b1011000000000000000000010000000,
31'b0000101000000000001010000100000,
31'b1100000000100000001010000000000,
31'b1100010000001000000000000000100,
31'b0011100000000000000010000100000,
31'b1000001000000000001000010000000,
31'b1001000000000000000010000000101,
31'b1100010000000000000000000000100,
31'b0010010000000001000000100000000,
31'b1100010000000100000000000000100,
31'b0011000010000000000100000000001,
31'b0000100000100000000010000001000,
31'b0000000000010000100000001001000,
31'b0000000010000000001000001000000,
31'b0000000000000001000010000000100,
31'b0000101010000000000101000000000,
31'b0010000001000100000000101000000,
31'b0000000010001000001000001000000,
31'b0010000001000000000000101000000,
31'b0000010000100001001000000000000,
31'b0000000000000000100000001001000,
31'b0000010000000000100010000000010,
31'b0000000000010001000010000000100,
31'b1000010000000000100000000010001,
31'b0010000000000001000000010000001,
31'b0001000110000000000100000000010,
31'b0010000001010000000000101000000,
31'b0000100000000000000010000001000,
31'b0000100000000010000010000001000,
31'b0000100000000100000010000001000,
31'b0000110000000000000000001000010,
31'b0000100000001000000010000001000,
31'b0100100000000000000001000010010,
31'b0000100001000000000001001000001,
31'b0011011000000001000000000000000,
31'b0000010000000001001000000000000,
31'b0000010000000011001000000000000,
31'b0000010000000101001000000000000,
31'b0000110000010000000000001000010,
31'b1000000000000000000000010101000,
31'b1010010000000000000100001000000,
31'b1000011100000000000000000000010,
31'b1010001000000000000000110000000,
31'b0000100010000000010000000100001,
31'b0010000000001100000000101000000,
31'b0000000011000000001000001000000,
31'b0010000000001000000000101000000,
31'b0000001000000000000000001101000,
31'b0010000000000100000000101000000,
31'b0000000000000000010110000000000,
31'b0010000000000000000000101000000,
31'b0101010000000000100001000000000,
31'b0000000100000001000001100000000,
31'b0001010000000000001100010000000,
31'b0010000100000000000000000001101,
31'b1100000000000000100010000001000,
31'b0010000001000001000000010000001,
31'b0001000000000000100000001010000,
31'b0010000000010000000000101000000,
31'b0000100001000000000010000001000,
31'b1001100000000000000000000000011,
31'b0000100001000100000010000001000,
31'b0011000000000000000000000100110,
31'b0000100001001000000010000001000,
31'b1100100000000000000000001001000,
31'b0000100000000000000001001000001,
31'b0010000000100000000000101000000,
31'b0100001100000000000000000001000,
31'b0100010000000000010000101000000,
31'b1000001010000000001000010000000,
31'b1001000000000000000000010110000,
31'b1100010010000000000000000000100,
31'b0011000000000100000100000000001,
31'b0011000000000010000100000000001,
31'b0011000000000000000100000000001,
31'b1011101000000000000000000000000,
31'b0010000000000000001100000000010,
31'b0001000000000011000001000000000,
31'b0001000000000001000001000000000,
31'b1000000000000001000000001000010,
31'b1000100000010100001000000000000,
31'b1000100000010010001000000000000,
31'b1000100000010000001000000000000,
31'b0100000011100000000000000001000,
31'b1000100000001100001000000000000,
31'b1010000100000000000001000000010,
31'b1000100000001000001000000000000,
31'b1000100000000110001000000000000,
31'b1000100000000100001000000000000,
31'b1000100000000010001000000000000,
31'b1000100000000000001000000000000,
31'b0111000000000010000000000100000,
31'b0111000000000000000000000100000,
31'b0101001000000000000000100001000,
31'b0100000001000000101000000000000,
31'b1000110000000000000010000000100,
31'b0111000000001000000000000100000,
31'b1000010010010000000000000000010,
31'b1000100000110000001000000000000,
31'b0100000011000000000000000001000,
31'b0111000000010000000000000100000,
31'b1000010010001000000000000000010,
31'b1000100000101000001000000000000,
31'b1000010010000100000000000000010,
31'b1000100000100100001000000000000,
31'b1000010010000000000000000000010,
31'b1000100000100000001000000000000,
31'b0100000010110000000000000001000,
31'b0100000000000001000010000000010,
31'b0100010000000001000000001001000,
31'b0100000000100000101000000000000,
31'b0000000010000000000100100000010,
31'b0100001000100000000000100010000,
31'b0010010010000000010000000001000,
31'b1100000000000001000000000010001,
31'b0100000010100000000000000001000,
31'b0100000010100010000000000001000,
31'b1010100010000000000000100000000,
31'b1000100001001000001000000000000,
31'b0100001000000000000111000000000,
31'b1000100001000100001000000000000,
31'b1000100001000010001000000000000,
31'b1000100001000000001000000000000,
31'b0100000010010000000000000001000,
31'b0000000000000000000101010000000,
31'b0100000000000010101000000000000,
31'b0100000000000000101000000000000,
31'b0100001000000010000000100010000,
31'b0100001000000000000000100010000,
31'b0110000000000000000000000111000,
31'b0100000000001000101000000000000,
31'b0100000010000000000000000001000,
31'b0100000010000010000000000001000,
31'b1000000100000000001000010000000,
31'b1000000010000000000001000000001,
31'b0100000010001000000000000001000,
31'b0100001000010000000000100010000,
31'b1000010011000000000000000000010,
31'b1000100001100000001000000000000,
31'b1110000000000000010000000000010,
31'b0011010000000000010000000010000,
31'b0001001000000000000010010010000,
31'b0001000010000001000001000000000,
31'b1000100000000000100000000001000,
31'b1000100000000010100000000001000,
31'b1000100000000100100000000001000,
31'b1000100010010000001000000000000,
31'b0100000001100000000000000001000,
31'b0101000100000001010000000000000,
31'b1010100001000000000000100000000,
31'b1000100010001000001000000000000,
31'b1000100000010000100000000001000,
31'b1000100010000100001000000000000,
31'b1000010000100000000000000000010,
31'b1000100010000000001000000000000,
31'b0100000001010000000000000001000,
31'b0111000010000000000000000100000,
31'b1000010000011000000000000000010,
31'b1000000001010000000001000000001,
31'b1000100000100000100000000001000,
31'b1000000000010000000010001001000,
31'b1000010000010000000000000000010,
31'b1000000000000001100000000000100,
31'b0100000001000000000000000001000,
31'b0100000001000010000000000001000,
31'b1000010000001000000000000000010,
31'b1000000001000000000001000000001,
31'b1000010000000100000000000000010,
31'b1000000000000000000010001001000,
31'b1000010000000000000000000000010,
31'b0101000000000000000000000010000,
31'b0100000000110000000000000001000,
31'b0100000010000001000010000000010,
31'b1010100000010000000000100000000,
31'b1001100000000000100000000010000,
31'b0000000000000000000100100000010,
31'b0000001000000000000010010001000,
31'b0010010000000000010000000001000,
31'b0010010000000010010000000001000,
31'b0100000000100000000000000001000,
31'b0100000000100010000000000001000,
31'b1010100000000000000000100000000,
31'b1000000000100000000001000000001,
31'b0100000000101000000000000001000,
31'b0100000000101010000000000001000,
31'b1010100000001000000000100000000,
31'b1000100011000000001000000000000,
31'b0100000000010000000000000001000,
31'b0100000000010010000000000001000,
31'b1000000000000000110100000000000,
31'b1000000000010000000001000000001,
31'b0100000000011000000000000001000,
31'b0100001010000000000000100010000,
31'b1000010001010000000000000000010,
31'b1000000001000001100000000000100,
31'b0100000000000000000000000001000,
31'b0100000000000010000000000001000,
31'b0100000000000100000000000001000,
31'b1000000000000000000001000000001,
31'b0100000000001000000000000001000,
31'b0100000000001010000000000001000,
31'b1000010001000000000000000000010,
31'b1000000000001000000001000000001,
31'b0000100000001000000101000000000,
31'b0011000000011000000000001000000,
31'b0000001000000000001000001000000,
31'b0001000100000001000001000000000,
31'b0000100000000000000101000000000,
31'b0011000000010000000000001000000,
31'b0000100000000100000101000000000,
31'b1010001000000001000100000000000,
31'b1010000000000100000001000000010,
31'b0011000000001000000000001000000,
31'b1010000000000000000001000000010,
31'b1010000000000010000001000000010,
31'b0011000000000010000000001000000,
31'b0011000000000000000000001000000,
31'b1010000000001000000001000000010,
31'b1000100100000000001000000000000,
31'b0000101010000000000010000001000,
31'b1100000001000000010000000000001,
31'b0000001000100000001000001000000,
31'b0101010000000000010000001000000,
31'b0000100000100000000101000000000,
31'b0010000000000000000100100000001,
31'b0000100001000000001010000100000,
31'b0011010010000001000000000000000,
31'b1100000000000001000000000100010,
31'b0011000000101000000000001000000,
31'b1000000001000000001000010000000,
31'b1000100000000000000000100000011,
31'b0011000000100010000000001000000,
31'b0011000000100000000000001000000,
31'b1000010110000000000000000000010,
31'b1010000010000000000000110000000,
31'b0000101000000000010000000100001,
31'b1100000000100000010000000000001,
31'b0000001001000000001000001000000,
31'b0100001000000001010000100000000,
31'b0000100001000000000101000000000,
31'b0011000001010000000000001000000,
31'b0000100001000100000101000000000,
31'b1100001000000000001010000000000,
31'b1111000000000000000010000000000,
31'b0011000001001000000000001000000,
31'b1000000000100000001000010000000,
31'b1010010000001000000000000000001,
31'b0110010000000000000001000001000,
31'b0011000001000000000000001000000,
31'b1010010000000010000000000000001,
31'b1010010000000000000000000000001,
31'b0000000010000000001100000000001,
31'b1100000000000000010000000000001,
31'b0000000000000000010001000001000,
31'b0100000100000000101000000000000,
31'b0000100001100000000101000000000,
31'b1100000000001000010000000000001,
31'b0000100000000000001010000100000,
31'b0100000100001000101000000000000,
31'b1000000000000100001000010000000,
31'b1100000000010000010000000000001,
31'b1000000000000000001000010000000,
31'b1000000000000010001000010000000,
31'b1100011000000000000000000000100,
31'b0011000001100000000000001000000,
31'b1000000000001000001000010000000,
31'b1010010000100000000000000000001,
31'b0000101000100000000010000001000,
31'b1100000000000000000010000101000,
31'b0000001010000000001000001000000,
31'b0001000000000000000000001110000,
31'b0000100010000000000101000000000,
31'b0101010000000000000001000100000,
31'b0000100010000100000101000000000,
31'b0011010000100001000000000000000,
31'b0101000000000011010000000000000,
31'b0101000000000001010000000000000,
31'b1010000010000000000001000000010,
31'b0101000000000101010000000000000,
31'b0101000001000000000100000000100,
31'b0100100000000000000000010001000,
31'b1000100000000000000001010000001,
31'b1010000000100000000000110000000,
31'b0000101000000000000010000001000,
31'b1000000001000000100000010001000,
31'b0000101000000100000010000001000,
31'b0011010000001001000000000000000,
31'b0000101000001000000010000001000,
31'b0011010000000101000000000000000,
31'b1001000000000000100000010010000,
31'b0011010000000001000000000000000,
31'b0100000101000000000000000001000,
31'b0101000000100001010000000000000,
31'b1000010100001000000000000000010,
31'b1010000000001000000000110000000,
31'b1000010100000100000000000000010,
31'b1010000000000100000000110000000,
31'b1000010100000000000000000000010,
31'b1010000000000000000000110000000,
31'b0000000000100000001100000000001,
31'b1000010000000000000000000110001,
31'b0000001011000000001000001000000,
31'b0010110000000000000000000010100,
31'b0000000000000000000000001101000,
31'b0010010000000000000100010000000,
31'b0000001000000000010110000000000,
31'b0010001000000000000000101000000,
31'b0100000100100000000000000001000,
31'b0101000001000001010000000000000,
31'b1010100100000000000000100000000,
31'b1000110000000000000000010000010,
31'b0101000000000000000100000000100,
31'b0101000000000010000100000000100,
31'b0101000000000100000100000000100,
31'b1010010010000000000000000000001,
31'b0000000000000000001100000000001,
31'b1000000000000000100000010001000,
31'b0000000010000000010001000001000,
31'b1000000100010000000001000000001,
31'b0000000000100000000000001101000,
31'b1010000000000001000000001000001,
31'b0000101000000000000001001000001,
31'b0011010001000001000000000000000,
31'b0100000100000000000000000001000,
31'b0100000100000010000000000001000,
31'b1000000010000000001000010000000,
31'b1000000100000000000001000000001,
31'b0100000100001000000000000001000,
31'b0100100000000000010000000010100,
31'b1000010101000000000000000000010,
31'b1010000001000000000000110000000,
31'b0010000000000000011000000100000,
31'b0110100000000000000000000010010,
31'b0001000001000000110000000000000,
31'b0001011000000001000001000000000,
31'b0100000100000000001001000010000,
31'b0100000000000000000010000100100,
31'b0001010000010000000100000000010,
31'b1100000000010000000100000010000,
31'b0010100000000001000000110000000,
31'b1100100000000000000000010000100,
31'b0001010000001000000100000000010,
31'b1100000000001000000100000010000,
31'b0011000000000000010000100001000,
31'b1100000000000100000100000010000,
31'b0001010000000000000100000000010,
31'b1100000000000000000100000010000,
31'b0010101010000000000100000000000,
31'b0000000100010000000010001000100,
31'b0101010000000000000000100001000,
31'b0000000100000001100000000001000,
31'b1001000001000000000000100000010,
31'b0000000001000000100000010000100,
31'b1100000000000000000011100000000,
31'b0010000100000000000000011000001,
31'b0000001000000000000000010100100,
31'b0000000100000000000010001000100,
31'b1100000000000001000000010001000,
31'b0010000001000000100010000000001,
31'b1100000101000000000000000000100,
31'b0010000101000001000000100000000,
31'b1000001010000000000000000000010,
31'b1100000000100000000100000010000,
31'b1000000000000000000000001100100,
31'b1001000010000000000001010000000,
31'b0001000000000000110000000000000,
31'b0001000000000010110000000000000,
31'b1001000000100000000000100000010,
31'b0000000010000000010000100100000,
31'b0001000000001000110000000000000,
31'b0001000000001010110000000000000,
31'b1101000000000000000100000001000,
31'b0010000000000100010000100010000,
31'b0001000000010000110000000000000,
31'b0010000000000000010000100010000,
31'b1100000100100000000000000000100,
31'b0010001000000000111000000000000,
31'b0001010001000000000100000000010,
31'b1100000001000000000100000010000,
31'b1001000000001000000000100000010,
31'b0000000000001000100000010000100,
31'b0001000000100000110000000000000,
31'b0000000000000000000001101000000,
31'b1001000000000000000000100000010,
31'b0000000000000000100000010000100,
31'b1001000000000100000000100000010,
31'b0000000000001000000001101000000,
31'b1100000100001000000000000000100,
31'b0010000100001001000000100000000,
31'b0011100000000000000100100000000,
31'b0010000000000000100010000000001,
31'b1100000100000000000000000000100,
31'b0010000100000001000000100000000,
31'b1100000100000100000000000000100,
31'b0010000100000101000000100000000,
31'b0010101000100000000100000000000,
31'b1110000000000000000100000100000,
31'b0001010000000000000010010010000,
31'b1100000000000000000010010000010,
31'b0100000000000010000000010010001,
31'b0100000000000000000000010010001,
31'b0000000001000000000000011000010,
31'b0100100000010000000000000100010,
31'b0000001000000000110000100000000,
31'b0001001000100000000001001000000,
31'b0000000100000000100010000000010,
31'b0110000000000000000010000010100,
31'b0000000000000100011000000010000,
31'b0100100000000100000000000100010,
31'b0000000000000000011000000010000,
31'b0100100000000000000000000100010,
31'b0010101000000000000100000000000,
31'b1011000000000000001000000000010,
31'b1000001000011000000000000000010,
31'b1000000000000001000101000000000,
31'b1001100100000000000001000000000,
31'b0100010000000000100000000101000,
31'b1000001000010000000000000000010,
31'b1000001000010010000000000000010,
31'b0000000100000001001000000000000,
31'b0001001000000000000001001000000,
31'b1000001000001000000000000000010,
31'b1000001000001010000000000000010,
31'b1000001000000100000000000000010,
31'b1010000100000000000100001000000,
31'b1000001000000000000000000000010,
31'b1000001000000010000000000000010,
31'b1001000000000010000001010000000,
31'b1001000000000000000001010000000,
31'b0001000010000000110000000000000,
31'b1001000000000100000001010000000,
31'b0000000000000100000000011000010,
31'b0000000000000000010000100100000,
31'b0000000000000000000000011000010,
31'b0000000000000100010000100100000,
31'b0101000100000000100001000000000,
31'b0001000000000000011000000001000,
31'b0001000100000000001100010000000,
31'b0010010000000000000000000001101,
31'b0000100000000011001000010000000,
31'b0000100000000001001000010000000,
31'b0000000001000000011000000010000,
31'b0100100001000000000000000100010,
31'b0100100100000000000000000010001,
31'b1001000000100000000001010000000,
31'b1000000000001000010001000000100,
31'b1000000000000000100000000100010,
31'b1001000010000000000000100000010,
31'b0000000010000000100000010000100,
31'b1000000000000000010001000000100,
31'b1000000000001000100000000100010,
31'b0100011000000000000000000001000,
31'b0100011000000010000000000001000,
31'b1000010000000001000000000100100,
31'b1000011000000000000001000000001,
31'b1100000110000000000000000000100,
31'b0010100000000000100100000100000,
31'b1000001001000000000000000000010,
31'b1000001001000010000000000000010,
31'b0000100000000000100000000000100,
31'b0000100000000010100000000000100,
31'b0000010000000000001000001000000,
31'b0000010000000010001000001000000,
31'b0100000000000000001001000010000,
31'b0100000100000000000010000100100,
31'b0000010000001000001000001000000,
31'b1010010000000001000100000000000,
31'b0000100000010000100000000000100,
31'b0000110000000001000000000000010,
31'b0000010000010000001000001000000,
31'b0000110000000101000000000000010,
31'b1100000001100000000000000000100,
31'b0011011000000000000000001000000,
31'b0001010100000000000100000000010,
31'b1100000100000000000100000010000,
31'b0000100000100000100000000000100,
31'b0000000000010000000010001000100,
31'b0000010000100000001000001000000,
31'b0000000000000001100000000001000,
31'b1100000001010000000000000000100,
31'b0010000001010001000000100000000,
31'b0010000000000010000000011000001,
31'b0010000000000000000000011000001,
31'b0000000010000001001000000000000,
31'b0000000000000000000010001000100,
31'b0000010000000000000000000001110,
31'b0000000000010001100000000001000,
31'b1100000001000000000000000000100,
31'b0010000001000001000000100000000,
31'b1100000001000100000000000000100,
31'b0010000001000101000000100000000,
31'b1001000000000000001000000000001,
31'b1001000000000010001000000000001,
31'b0001000100000000110000000000000,
31'b0101000000000000001001000001000,
31'b1100000000110000000000000000100,
31'b0010001010000000000100010000000,
31'b0001000100001000110000000000000,
31'b1100010000000000001010000000000,
31'b1100000000101000000000000000100,
31'b0010001000000000000010000010010,
31'b0001000100010000110000000000000,
31'b1101000000000000010000010000000,
31'b1100000000100000000000000000100,
31'b0010000000100001000000100000000,
31'b1100000000100100000000000000100,
31'b1010001000000000000000000000001,
31'b1100000000011000000000000000100,
31'b0010000000011001000000100000000,
31'b0001001000000001001000100000000,
31'b0000000100000000000001101000000,
31'b1100000000010000000000000000100,
31'b0010000000010001000000100000000,
31'b1100000000010100000000000000100,
31'b0010000001000000000000011000001,
31'b1100000000001000000000000000100,
31'b0010000000001001000000100000000,
31'b1100000000001100000000000000100,
31'b0010000100000000100010000000001,
31'b1100000000000000000000000000100,
31'b0010000000000001000000100000000,
31'b1100000000000100000000000000100,
31'b0010000000000101000000100000000,
31'b0000100010000000100000000000100,
31'b0000100010000010100000000000100,
31'b0000010010000000001000001000000,
31'b0000100000100000000000001000010,
31'b1001100000100000000001000000000,
31'b1011000000000000000000100000001,
31'b0000010010001000001000001000000,
31'b0011001000100001000000000000000,
31'b0000000000100001001000000000000,
31'b0000010000000000100000001001000,
31'b0000000000000000100010000000010,
31'b0000100000000000001000000001100,
31'b1000000000000000100000000010001,
31'b1010000000100000000100001000000,
31'b0000000100000000011000000010000,
31'b0100100100000000000000000100010,
31'b0000000000010001001000000000000,
31'b0000100000000100000000001000010,
31'b0000100000000010000000001000010,
31'b0000100000000000000000001000010,
31'b1001100000000000000001000000000,
31'b1010000000010000000100001000000,
31'b1001100000000100000001000000000,
31'b0011001000000001000000000000000,
31'b0000000000000001001000000000000,
31'b0000000000000011001000000000000,
31'b0000000000000101001000000000000,
31'b0000100000010000000000001000010,
31'b0000000000001001001000000000000,
31'b1010000000000000000100001000000,
31'b1000001100000000000000000000010,
31'b1010000000000100000100001000000,
31'b1001000010000000001000000000001,
31'b1001000100000000000001010000000,
31'b0001000110000000110000000000000,
31'b0010101000000000000000000010100,
31'b0010001000000010000100010000000,
31'b0010001000000000000100010000000,
31'b0000010000000000010110000000000,
31'b0010010000000000000000101000000,
31'b0101000000000000100001000000000,
31'b0101000000000010100001000000000,
31'b0001000000000000001100010000000,
31'b1001000000000000100000000001001,
31'b1100000010100000000000000000100,
31'b0010001000010000000100010000000,
31'b0001010000000000100000001010000,
31'b1100000000000000100000001000010,
31'b0100100000000000000000000010001,
31'b0100100000000010000000000010001,
31'b0100100000000100000000000010001,
31'b0000100001000000000000001000010,
31'b1100000010010000000000000000100,
31'b0010001000100000000100010000000,
31'b1100100000000000000010000000010,
31'b0011001001000001000000000000000,
31'b0000000001000001001000000000000,
31'b0100000000000000010000101000000,
31'b0100000000000000000000010100010,
31'b0100000000000100010000101000000,
31'b1100000010000000000000000000100,
31'b0010000010000001000000100000000,
31'b1100000010000100000000000000100,
31'b0011010000000000000100000000001,
31'b0010100010100000000100000000000,
31'b0011000010000000010000000010000,
31'b0100000100000000100001100000000,
31'b0001010000000001000001000000000,
31'b1000100000100000000010000000100,
31'b1000000000010000100000001000100,
31'b1000000010110000000000000000010,
31'b1000000000000001000010000001000,
31'b0000000010000000110000100000000,
31'b1000000000001000100000001000100,
31'b1000000010101000000000000000010,
31'b1000000000000000000001110000000,
31'b1000000010100100000000000000010,
31'b1000000000000000100000001000100,
31'b1000000010100000000000000000010,
31'b0001000000000000010000000100000,
31'b0010100010000000000100000000000,
31'b0111010000000000000000000100000,
31'b1000000010011000000000000000010,
31'b0101000100000000010000001000000,
31'b1000100000000000000010000000100,
31'b1000100000000010000010000000100,
31'b1000000010010000000000000000010,
31'b1000000010010010000000000000010,
31'b0000000000000000000000010100100,
31'b0001000010000000000001001000000,
31'b1000000010001000000000000000010,
31'b1000000010001010000000000000010,
31'b1000000010000100000000000000010,
31'b1000000010000110000000000000010,
31'b1000000010000000000000000000010,
31'b1000000010000010000000000000010,
31'b1001000000000001000010000010000,
31'b1000000100000000000010010000100,
31'b0100000000000001000000001001000,
31'b0100010000100000101000000000000,
31'b0010000010000100010000000001000,
31'b0010000110000000000100010000000,
31'b0010000010000000010000000001000,
31'b1010000100010000000000000000001,
31'b0100000000000000100010000000100,
31'b0100100000000000001000000001010,
31'b0100000000010001000000001001000,
31'b1010000100001000000000000000001,
31'b0110000100000000000001000001000,
31'b0010000000000000111000000000000,
31'b1010000100000010000000000000001,
31'b1010000100000000000000000000001,
31'b0100100000000010000000001000100,
31'b0100100000000000000000001000100,
31'b0100010000000010101000000000000,
31'b0100010000000000101000000000000,
31'b1001001000000000000000100000010,
31'b0000100000000000001100100000000,
31'b1001000100000000010010000000000,
31'b0100010000001000101000000000000,
31'b0100010010000000000000000001000,
31'b0100100000010000000000001000100,
31'b1000010100000000001000010000000,
31'b1010000000000000001000100000010,
31'b1100001100000000000000000000100,
31'b0010001100000001000000100000000,
31'b1000000011000000000000000000010,
31'b1010000100100000000000000000001,
31'b0010100000100000000100000000000,
31'b0011000000000000010000000010000,
31'b1100000000000000000100100001000,
31'b0011000000000100010000000010000,
31'b1000110000000000100000000001000,
31'b0101000100000000000001000100000,
31'b1000000000110000000000000000010,
31'b1000000010000001000010000001000,
31'b0000000000000000110000100000000,
31'b0001000000100000000001001000000,
31'b1000000000101000000000000000010,
31'b1000000010000000000001110000000,
31'b1000000000100100000000000000010,
31'b1000000010000000100000001000100,
31'b1000000000100000000000000000010,
31'b1000000000100010000000000000010,
31'b0010100000000000000100000000000,
31'b0010100000000010000100000000000,
31'b1000000000011000000000000000010,
31'b1000001000000001000101000000000,
31'b1000000000010100000000000000010,
31'b1000100000000001001000001000000,
31'b1000000000010000000000000000010,
31'b1000000000010010000000000000010,
31'b0000000000000000000010000010001,
31'b0001000000000000000001001000000,
31'b1000000000001000000000000000010,
31'b1000000000001010000000000000010,
31'b1000000000000100000000000000010,
31'b1000000000000110000000000000010,
31'b1000000000000000000000000000010,
31'b1000000000000010000000000000010,
31'b0100100000000100100000000000010,
31'b1001001000000000000001010000000,
31'b0100100000000000100000000000010,
31'b0100100000000010100000000000010,
31'b0010000000000100010000000001000,
31'b0010000100000000000100010000000,
31'b0010000000000000010000000001000,
31'b0010000000000010010000000001000,
31'b0100010000100000000000000001000,
31'b0100010000100010000000000001000,
31'b1010110000000000000000100000000,
31'b1000100100000000000000010000010,
31'b1110000000000000100100000000000,
31'b0010000100010000000100010000000,
31'b1000000001100000000000000000010,
31'b1010000110000000000000000000001,
31'b0100010000010000000000000001000,
31'b0100100010000000000000001000100,
31'b1000010000000000110100000000000,
31'b1000010000010000000001000000001,
31'b1100100000000000010000100000000,
31'b0010100000000001010000000000100,
31'b1000000001010000000000000000010,
31'b1000000001010010000000000000010,
31'b0100010000000000000000000001000,
31'b0100010000000010000000000001000,
31'b1000000001001000000000000000010,
31'b1000010000000000000001000000001,
31'b1000000001000100000000000000010,
31'b1100000000000000000000001010001,
31'b1000000001000000000000000000010,
31'b1000000001000010000000000000010,
31'b0000101000000000100000000000100,
31'b1000000001000000000010010000100,
31'b0100000000000000100001100000000,
31'b0101000000100000010000001000000,
31'b0100000000000000000000011000100,
31'b0101000010000000000001000100000,
31'b0100000000001000100001100000000,
31'b1010000001010000000000000000001,
31'b0000101000010000100000000000100,
31'b0011010000001000000000001000000,
31'b1010010000000000000001000000010,
31'b1010000001001000000000000000001,
31'b0110000001000000000001000001000,
31'b0011010000000000000000001000000,
31'b1010000001000010000000000000001,
31'b1010000001000000000000000000001,
31'b0010100110000000000100000000000,
31'b1100000000000000100000000100100,
31'b0101000000000010010000001000000,
31'b0101000000000000010000001000000,
31'b1100000000000000010001000000010,
31'b0011000010000101000000000000000,
31'b1001000001000000010010000000000,
31'b0011000010000001000000000000000,
31'b0000001010000001001000000000000,
31'b0001000000000001000000000110000,
31'b1000010001000000001000010000000,
31'b0101000000010000010000001000000,
31'b1100001001000000000000000000100,
31'b0011010000100000000000001000000,
31'b1000000110000000000000000000010,
31'b1010000001100000000000000000001,
31'b1001001000000000001000000000001,
31'b1000000000000000000010010000100,
31'b0100000100000001000000001001000,
31'b1010000000011000000000000000001,
31'b0110000000010000000001000001000,
31'b0010000010000000000100010000000,
31'b1010000000010010000000000000001,
31'b1010000000010000000000000000001,
31'b0110000000001000000001000001000,
31'b0010000000000000000010000010010,
31'b1010000000001010000000000000001,
31'b1010000000001000000000000000001,
31'b0110000000000000000001000001000,
31'b0000100000000000000000000100100,
31'b1010000000000010000000000000001,
31'b1010000000000000000000000000001,
31'b0010000010000001000000000011000,
31'b1100010000000000010000000000001,
31'b0001000000000001001000100000000,
31'b0101000001000000010000001000000,
31'b1100001000010000000000000000100,
31'b0010001000010001000000100000000,
31'b1001000000000000010010000000000,
31'b1010000000110000000000000000001,
31'b1100001000001000000000000000100,
31'b0010001000001001000000100000000,
31'b1000010000000000001000010000000,
31'b1010000000101000000000000000001,
31'b1100001000000000000000000000100,
31'b0010001000000001000000100000000,
31'b0000000000000001000000000101000,
31'b1010000000100000000000000000001,
31'b0010100100100000000100000000000,
31'b1100000000000000010000110000000,
31'b1100000000000000000000001100010,
31'b0011000000101001000000000000000,
31'b0101000000000010000001000100000,
31'b0101000000000000000001000100000,
31'b1001000000000000000000000101001,
31'b0011000000100001000000000000000,
31'b0000001000100001001000000000000,
31'b0101010000000001010000000000000,
31'b1000000000000000001000100000001,
31'b1000100001000000000000010000010,
31'b1000001000000000100000000010001,
31'b0101000000010000000001000100000,
31'b1000000100100000000000000000010,
31'b1010000011000000000000000000001,
31'b0010100100000000000100000000000,
31'b0011000000001101000000000000000,
31'b1001000000000000001100001000000,
31'b0011000000001001000000000000000,
31'b1001101000000000000001000000000,
31'b0011000000000101000000000000000,
31'b1000000100010000000000000000010,
31'b0011000000000001000000000000000,
31'b0000001000000001001000000000000,
31'b0001000100000000000001001000000,
31'b1000000100001000000000000000010,
31'b1010100000000000001001000000000,
31'b1000000100000100000000000000010,
31'b1010001000000000000100001000000,
31'b1000000100000000000000000000010,
31'b1000000100000010000000000000010,
31'b1000000000000010000000000110001,
31'b1000000000000000000000000110001,
31'b0100100100000000100000000000010,
31'b0010100000000000000000000010100,
31'b0010000000000010000100010000000,
31'b0010000000000000000100010000000,
31'b0010000100000000010000000001000,
31'b0000000000000000000010000100010,
31'b0101001000000000100001000000000,
31'b1000100000000100000000010000010,
31'b1000100000000010000000010000010,
31'b1000100000000000000000010000010,
31'b0110000010000000000001000001000,
31'b0010000000010000000100010000000,
31'b1010000010000010000000000000001,
31'b1010000010000000000000000000001,
31'b0010000000000001000000000011000,
31'b1000010000000000100000010001000,
31'b0011000000000000010100000000100,
31'b0011000001001001000000000000000,
31'b0010000000100010000100010000000,
31'b0010000000100000000100010000000,
31'b1001000010000000010010000000000,
31'b0011000001000001000000000000000,
31'b0100010100000000000000000001000,
31'b0100010100000010000000000001000,
31'b1000010010000000001000010000000,
31'b1000100000100000000000010000010,
31'b1100001010000000000000000000100,
31'b0010001010000001000000100000000,
31'b1000000101000000000000000000010,
31'b1010000010100000000000000000001,
31'b1100000000000000000000000000000,
31'b1100000000000010000000000000000,
31'b1100000000000100000000000000000,
31'b0000000000000000000001000001001,
31'b1100000000001000000000000000000,
31'b0000000001000000000010001000000,
31'b1100000000001100000000000000000,
31'b0000000001000100000010001000000,
31'b1100000000010000000000000000000,
31'b0000000100000000100000010000000,
31'b1100000000010100000000000000000,
31'b0000000100000100100000010000000,
31'b1100000000011000000000000000000,
31'b0000000100001000100000010000000,
31'b1100000000011100000000000000000,
31'b0000000100001100100000010000000,
31'b1100000000100000000000000000000,
31'b0000101000000000000000000100000,
31'b1100000000100100000000000000000,
31'b0000101000000100000000000100000,
31'b1100000000101000000000000000000,
31'b0000101000001000000000000100000,
31'b1100000000101100000000000000000,
31'b0000101000001100000000000100000,
31'b1100000000110000000000000000000,
31'b0000101000010000000000000100000,
31'b1100000000110100000000000000000,
31'b0001100000000000100000000011000,
31'b0000100001000000100000000000000,
31'b1000001000000000000010010000000,
31'b1010010000000000010000000000000,
31'b1010010000000010010000000000000,
31'b1100000001000000000000000000000,
31'b0000000000001000000010001000000,
31'b1100000001000100000000000000000,
31'b0000000001000000000001000001001,
31'b0000000000000010000010001000000,
31'b0000000000000000000010001000000,
31'b0000010000000000000000000001010,
31'b0000000000000100000010001000000,
31'b1100000001010000000000000000000,
31'b0000000101000000100000010000000,
31'b1100000001010100000000000000000,
31'b0010000100000001000011000000000,
31'b0000100000100000100000000000000,
31'b0000000000010000000010001000000,
31'b0000100000100100100000000000000,
31'b0000000000010100000010001000000,
31'b1100000001100000000000000000000,
31'b0000101001000000000000000100000,
31'b1100000001100100000000000000000,
31'b0000101001000100000000000100000,
31'b0000100000010000100000000000000,
31'b0000000000100000000010001000000,
31'b0000100000010100100000000000000,
31'b0000100010000000001000000001000,
31'b0000100000001000100000000000000,
31'b0100000100000000000010000100000,
31'b0100010000000000000100100000000,
31'b0100010000000010000100100000000,
31'b0000100000000000100000000000000,
31'b0000100000000010100000000000000,
31'b0000100000000100100000000000000,
31'b0000100000000110100000000000000,
31'b1100000010000000000000000000000,
31'b0000000000000000011100000000000,
31'b1100000010000100000000000000000,
31'b0000000010000000000001000001001,
31'b1100000010001000000000000000000,
31'b0000000011000000000010001000000,
31'b1100000010001100000000000000000,
31'b0000101000000000010001001000000,
31'b1100000010010000000000000000000,
31'b0000000110000000100000010000000,
31'b1000000100000000010001000000000,
31'b1100000000000000101000000001000,
31'b1100000010011000000000000000000,
31'b0001010000000000000110010000000,
31'b1110000000000000000000000110000,
31'b0011010000000000000000000100010,
31'b1100000010100000000000000000000,
31'b0000101010000000000000000100000,
31'b1100000010100100000000000000000,
31'b0000101010000100000000000100000,
31'b1100000010101000000000000000000,
31'b0000101010001000000000000100000,
31'b0001101000000000100000100000000,
31'b0000100001000000001000000001000,
31'b1100000010110000000000000000000,
31'b0010100000000000101000100000000,
31'b1100010000000001000000001000000,
31'b0010101000001000000000000010000,
31'b1000000000000001000001000010000,
31'b1000001010000000000010010000000,
31'b1010010010000000010000000000000,
31'b0010101000000000000000000010000,
31'b1100000011000000000000000000000,
31'b0000000010001000000010001000000,
31'b1100000011000100000000000000000,
31'b0000100000101000001000000001000,
31'b0000000000000001001000000000100,
31'b0000000010000000000010001000000,
31'b0000010010000000000000000001010,
31'b0000100000100000001000000001000,
31'b1100000011010000000000000000000,
31'b0000010100000000010010000010000,
31'b1101001000000000000000100000000,
31'b0011001000000001000000000000100,
31'b0000100010100000100000000000000,
31'b0000010000000000101000000000010,
31'b0000100010100100100000000000000,
31'b0000100000000000000000001000110,
31'b1100000011100000000000000000000,
31'b0000101011000000000000000100000,
31'b0010100000000000100000000110000,
31'b0000100000001000001000000001000,
31'b0000100010010000100000000000000,
31'b0000100000000100001000000001000,
31'b0000100000000010001000000001000,
31'b0000100000000000001000000001000,
31'b0101000000000001000000000000001,
31'b0101000000000011000000000000001,
31'b0101000000000101000000000000001,
31'b0001100000000000000000100100000,
31'b0000100010000000100000000000000,
31'b0000100010000010100000000000000,
31'b0000100010000100100000000000000,
31'b0000010000000001000010000000000,
31'b1100000100000000000000000000000,
31'b0000000000010000100000010000000,
31'b1100000100000100000000000000000,
31'b0000000100000000000001000001001,
31'b1100000100001000000000000000000,
31'b0000000101000000000010001000000,
31'b1100000100001100000000000000000,
31'b0010000001000000000000110001000,
31'b0000000000000010100000010000000,
31'b0000000000000000100000010000000,
31'b1000000010000000010001000000000,
31'b0000000000000100100000010000000,
31'b1000000000100000000000001100000,
31'b0000000000001000100000010000000,
31'b1000000010001000010001000000000,
31'b0000000000001100100000010000000,
31'b1100000100100000000000000000000,
31'b0000101100000000000000000100000,
31'b1100000100100100000000000000000,
31'b0001011000000000100000000000001,
31'b1000000000010000000000001100000,
31'b1100100001000000000000010000000,
31'b1100000000000001010000000010000,
31'b0010010010000000000000000001001,
31'b1000000000001000000000001100000,
31'b0000000000100000100000010000000,
31'b1000000010100000010001000000000,
31'b0001000000000000000001000100010,
31'b1000000000000000000000001100000,
31'b1000000000000010000000001100000,
31'b1000000000000100000000001100000,
31'b1000000000000110000000001100000,
31'b1100000101000000000000000000000,
31'b0000000100001000000010001000000,
31'b1100000101000100000000000000000,
31'b0010000000010001000011000000000,
31'b0000001000000000000000010100000,
31'b0000000100000000000010001000000,
31'b0000010100000000000000000001010,
31'b0010000000000000000000110001000,
31'b1000101000000000000010000000000,
31'b0000000001000000100000010000000,
31'b1000101000000100000010000000000,
31'b0010000000000001000011000000000,
31'b0000100100100000100000000000000,
31'b0000000100010000000010001000000,
31'b0001010000100000000000000100001,
31'b0010000000010000000000110001000,
31'b1100000101100000000000000000000,
31'b1000001000000000100000001000000,
31'b0010000010000000000001000001010,
31'b1100000000000000000100000010100,
31'b0000100100010000100000000000000,
31'b1100100000000000000000010000000,
31'b0001010000010000000000000100001,
31'b1100100000000100000000010000000,
31'b0100000000000010000010000100000,
31'b0100000000000000000010000100000,
31'b0100010100000000000100100000000,
31'b0100000000000100000010000100000,
31'b0000100100000000100000000000000,
31'b0100000000001000000010000100000,
31'b0001010000000000000000000100001,
31'b0100100010000000000100000000001,
31'b1100000110000000000000000000000,
31'b0000000100000000011100000000000,
31'b0000000000000000001000010001000,
31'b1000000000000000100100000000001,
31'b1100000110001000000000000000000,
31'b0001000001000000001000010010000,
31'b1000010000000001000000000100000,
31'b1000010000000011000000000100000,
31'b1000000000000100010001000000000,
31'b0000000010000000100000010000000,
31'b1000000000000000010001000000000,
31'b1000000000000010010001000000000,
31'b1000000010100000000000001100000,
31'b0001000000000000010000001000010,
31'b1000000000001000010001000000000,
31'b1000000000001010010001000000000,
31'b1100000110100000000000000000000,
31'b0000101110000000000000000100000,
31'b1010000000000000000000001010000,
31'b1010000000000010000000001010000,
31'b1110010000000000000001000000000,
31'b0011000000000000000001000010010,
31'b1010000000001000000000001010000,
31'b0010010000000000000000000001001,
31'b1000000010001000000000001100000,
31'b0000000010100000100000010000000,
31'b1000000000100000010001000000000,
31'b1001000000000000100000101000000,
31'b1000000010000000000000001100000,
31'b1001000000000000000001010000100,
31'b1000000010000100000000001100000,
31'b0100100001000000000100000000001,
31'b1100000111000000000000000000000,
31'b0001010000000000100100001000000,
31'b1000001000000000000000000000110,
31'b1000001000000010000000000000110,
31'b0000001010000000000000010100000,
31'b0001000000000000001000010010000,
31'b1000010001000001000000000100000,
31'b0110000000100000000010000010000,
31'b1000101010000000000010000000000,
31'b0000010000000000010010000010000,
31'b1000000001000000010001000000000,
31'b1000011000000001100000000000000,
31'b0010101000000000000100000000100,
31'b0001000001000000010000001000010,
31'b1000001000000000000100000100001,
31'b1000010000000000010000000000011,
31'b0011010000000000000000000010001,
31'b1110000000000000000000000000011,
31'b0010000000000000000001000001010,
31'b0110000000001000000010000010000,
31'b0000100110010000100000000000000,
31'b1100100010000000000000010000000,
31'b0110000000000010000010000010000,
31'b0110000000000000000010000010000,
31'b0101000100000001000000000000001,
31'b0100000010000000000010000100000,
31'b1000001000000000001000001001000,
31'b0100100000001000000100000000001,
31'b0000100110000000100000000000000,
31'b0100100000000100000100000000001,
31'b0101000000000000100010100000000,
31'b0100100000000000000100000000001,
31'b1100001000000000000000000000000,
31'b0000100000100000000000000100000,
31'b1100001000000100000000000000000,
31'b0000100000100100000000000100000,
31'b1100001000001000000000000000000,
31'b0000100000101000000000000100000,
31'b1100001000001100000000000000000,
31'b0000100010000000010001001000000,
31'b1100001000010000000000000000000,
31'b0000100000110000000000000100000,
31'b1100001000010100000000000000000,
31'b0000110100000000000001000010000,
31'b1100001000011000000000000000000,
31'b1000000000100000000010010000000,
31'b0011000010000000010100000000000,
31'b1111000000000000001000000000000,
31'b0000100000000010000000000100000,
31'b0000100000000000000000000100000,
31'b0100000000000001000000100000001,
31'b0000100000000100000000000100000,
31'b0100000100000000100010000000000,
31'b0000100000001000000000000100000,
31'b0100000100000100100010000000000,
31'b0000100000001100000000000100000,
31'b0100000001000000000000011000000,
31'b0000100000010000000000000100000,
31'b0100000001000100000000011000000,
31'b0000100000010100000000000100000,
31'b1000000000000010000010010000000,
31'b1000000000000000000010010000000,
31'b1010011000000000010000000000000,
31'b1000000000000100000010010000000,
31'b1100001001000000000000000000000,
31'b0000100001100000000000000100000,
31'b1100001001000100000000000000000,
31'b0000100001100100000000000100000,
31'b0000000100000000000000010100000,
31'b0000001000000000000010001000000,
31'b0000011000000000000000000001010,
31'b0000001000000100000010001000000,
31'b1000100100000000000010000000000,
31'b1100000000001000100000000100000,
31'b1101000010000000000000100000000,
31'b0011000010000001000000000000100,
31'b0000101000100000100000000000000,
31'b1100000000000000100000000100000,
31'b0000101000100100100000000000000,
31'b1100000000000100100000000100000,
31'b0100000000010000000000011000000,
31'b0000100001000000000000000100000,
31'b0100000001000001000000100000001,
31'b0000100001000100000000000100000,
31'b0000101000010000100000000000000,
31'b0000100001001000000000000100000,
31'b0001100000000000000000000111000,
31'b0000101010000000001000000001000,
31'b0100000000000000000000011000000,
31'b0100000000000010000000011000000,
31'b0100000000000100000000011000000,
31'b0100000000000110000000011000000,
31'b0000101000000000100000000000000,
31'b1000000001000000000010010000000,
31'b0000101000000100100000000000000,
31'b1010000000000001100001000000000,
31'b1100001010000000000000000000000,
31'b0000100010100000000000000100000,
31'b1100001010000100000000000000000,
31'b0000100010100100000000000100000,
31'b1100001010001000000000000000000,
31'b0000100010101000000000000100000,
31'b0011000000010000010100000000000,
31'b0000100000000000010001001000000,
31'b1100001010010000000000000000000,
31'b0010100100000001010000000000000,
31'b1101000001000000000000100000000,
31'b0011000001000001000000000000100,
31'b0011000000000100010100000000000,
31'b1100000000000000000000100011000,
31'b0011000000000000010100000000000,
31'b0010100000100000000000000010000,
31'b0101010000000000000100000000000,
31'b0000100010000000000000000100000,
31'b0101010000000100000100000000000,
31'b0000100010000100000000000100000,
31'b0101010000001000000100000000000,
31'b0000100010001000000000000100000,
31'b0001100000000000100000100000000,
31'b0000000000000000000110000000001,
31'b0101010000010000000100000000000,
31'b0010000000000000000100010000100,
31'b0010100000001010000000000010000,
31'b0010100000001000000000000010000,
31'b1000001000000001000001000010000,
31'b1000000010000000000010010000000,
31'b0010100000000010000000000010000,
31'b0010100000000000000000000010000,
31'b1100001011000000000000000000000,
31'b0000100011100000000000000100000,
31'b1000000100000000000000000000110,
31'b1110000000000000100000000010000,
31'b0000001000000001001000000000100,
31'b0000001010000000000010001000000,
31'b1100000000000000001000000101000,
31'b0000101000100000001000000001000,
31'b1101000000000100000000100000000,
31'b0011000000000101000000000000100,
31'b1101000000000000000000100000000,
31'b0011000000000001000000000000100,
31'b0010100100000000000100000000100,
31'b1100000010000000100000000100000,
31'b1101000000001000000000100000000,
31'b0011000000001001000000000000100,
31'b0101010001000000000100000000000,
31'b0000100011000000000000000100000,
31'b1100000000000000000100001000001,
31'b0000101000001000001000000001000,
31'b0010100000000000001000100100000,
31'b0000101000000100001000000001000,
31'b1001000000000000000100000001010,
31'b0000101000000000001000000001000,
31'b0100000010000000000000011000000,
31'b0101000000000000000001000100100,
31'b1101000000100000000000100000000,
31'b0011000000100001000000000000100,
31'b0010000000000001010000010000000,
31'b1000010000000000110000000010000,
31'b0010100001000010000000000010000,
31'b0010100001000000000000000010000,
31'b1100001100000000000000000000000,
31'b0000100100100000000000000100000,
31'b1100001100000100000000000000000,
31'b0001010000100000100000000000001,
31'b0000000001000000000000010100000,
31'b0100100000010000000000001000000,
31'b0100000000000001001000000000010,
31'b0100100000010100000000001000000,
31'b1000100001000000000010000000000,
31'b0000001000000000100000010000000,
31'b1000100001000100000010000000000,
31'b0000110000000000000001000010000,
31'b0100100000000010000000001000000,
31'b0100100000000000000000001000000,
31'b0100100000000110000000001000000,
31'b0100100000000100000000001000000,
31'b0100000000001000100010000000000,
31'b0000100100000000000000000100000,
31'b0100000100000001000000100000001,
31'b0001010000000000100000000000001,
31'b0100000000000000100010000000000,
31'b0100000000000010100010000000000,
31'b0100000000000100100010000000000,
31'b0100110010000001000000000000000,
31'b1000100001100000000010000000000,
31'b0000100100010000000000000100000,
31'b0010010000000000000000100010001,
31'b0001010000010000100000000000001,
31'b1000001000000000000000001100000,
31'b1000000100000000000010010000000,
31'b1000001000000100000000001100000,
31'b1010000000000000000000101001000,
31'b0000000000001000000000010100000,
31'b1000000000100000100000001000000,
31'b1000000010000000000000000000110,
31'b1000000010000010000000000000110,
31'b0000000000000000000000010100000,
31'b0000000000000010000000010100000,
31'b0000000000000100000000010100000,
31'b0000000000000110000000010100000,
31'b1000100000000000000010000000000,
31'b1000100000000010000010000000000,
31'b1000100000000100000010000000000,
31'b1000100000000110000010000000000,
31'b0000000000010000000000010100000,
31'b0100100001000000000000001000000,
31'b0000100000000000000000000010011,
31'b0100100001000100000000001000000,
31'b1000000000000010100000001000000,
31'b1000000000000000100000001000000,
31'b1000000010100000000000000000110,
31'b1000000000000100100000001000000,
31'b0000000000100000000000010100000,
31'b1000000000001000100000001000000,
31'b0001000000000000100001000000010,
31'b1000000000001100100000001000000,
31'b1000100000100000000010000000000,
31'b1000000000010000100000001000000,
31'b1000100000100100000010000000000,
31'b1000000000010100100000001000000,
31'b0000101100000000100000000000000,
31'b1000000101000000000010010000000,
31'b0001011000000000000000000100001,
31'b0010000010000001000100000001000,
31'b1100001110000000000000000000000,
31'b0010100000010001010000000000000,
31'b1000000001000000000000000000110,
31'b1000001000000000100100000000001,
31'b0100010000000000000000000001100,
31'b0100100010010000000000001000000,
31'b1000011000000001000000000100000,
31'b1000010000000000000001000000101,
31'b1000100011000000000010000000000,
31'b0010100000000001010000000000000,
31'b1000001000000000010001000000000,
31'b1000010001000001100000000000000,
31'b0100100010000010000000001000000,
31'b0100100010000000000000001000000,
31'b1000001000001000010001000000000,
31'b0100100010000100000000001000000,
31'b0101010100000000000100000000000,
31'b0000100110000000000000000100000,
31'b1010001000000000000000001010000,
31'b0101000000000000000010100100000,
31'b0100000010000000100010000000000,
31'b0100110000000101000000000000000,
31'b0100110000000011000000000000000,
31'b0100110000000001000000000000000,
31'b0011000000000001000100000010000,
31'b0010100000100001010000000000000,
31'b0010000000000000010000000001100,
31'b0100100000000000010001000100000,
31'b1000001010000000000000001100000,
31'b1001000000000000001000001010000,
31'b0100100000000000100000000000110,
31'b0100000000000000001010000001000,
31'b1000000000000100000000000000110,
31'b1000000010100000100000001000000,
31'b1000000000000000000000000000110,
31'b1000000000000010000000000000110,
31'b0000000010000000000000010100000,
31'b0001000000000000000001001000100,
31'b1000000000001000000000000000110,
31'b1000000000001010000000000000110,
31'b1000100010000000000010000000000,
31'b1000100010000010000010000000000,
31'b0010000000000000000000010010000,
31'b1000010000000001100000000000000,
31'b0010100000000000000100000000100,
31'b0100100011000000000000001000000,
31'b1000000000000000000100000100001,
31'b1000010000001001100000000000000,
31'b1000000010000010100000001000000,
31'b1000000010000000100000001000000,
31'b1000000000100000000000000000110,
31'b1000000010000100100000001000000,
31'b0000000010100000000000010100000,
31'b1001000000000000010000010000010,
31'b1001000000000000000000101100000,
31'b0110001000000000000010000010000,
31'b1000100010100000000010000000000,
31'b1000010000000000001010000000010,
31'b1000000000000000001000001001000,
31'b1000010000100001100000000000000,
31'b0010100000100000000100000000100,
31'b0011000000000000010000000010100,
31'b1000000000100000000100000100001,
31'b0010000000000001000100000001000,
31'b1100010000000000000000000000000,
31'b0001000000000000000000000010010,
31'b1100010000000100000000000000000,
31'b0001000000000100000000000010010,
31'b1100010000001000000000000000000,
31'b0001000000001000000000000010010,
31'b0000000001000000000000000001010,
31'b1001000000000000000010000000001,
31'b1100010000010000000000000000000,
31'b0001000000010000000000000010010,
31'b1100010000010100000000000000000,
31'b0001100000000000000000010100001,
31'b1100010000011000000000000000000,
31'b0001000010000000000110010000000,
31'b1010000000100000010000000000000,
31'b1010000000100010010000000000000,
31'b1100010000100000000000000000000,
31'b0001000000100000000000000010010,
31'b1100010000100100000000000000000,
31'b0001001100000000100000000000001,
31'b1100010000101000000000000000000,
31'b0001001000000001000010100000000,
31'b1010000000010000010000000000000,
31'b1010000000010010010000000000000,
31'b1100010000110000000000000000000,
31'b0001001000000000000001010001000,
31'b1010000000001000010000000000000,
31'b1100000000000000001010000000100,
31'b1010000000000100010000000000000,
31'b1010000000000110010000000000000,
31'b1010000000000000010000000000000,
31'b1010000000000010010000000000000,
31'b1100010001000000000000000000000,
31'b0001000001000000000000000010010,
31'b0000000000001000000000000001010,
31'b0100000000000000000011000010000,
31'b0000000000000100000000000001010,
31'b0000010000000000000010001000000,
31'b0000000000000000000000000001010,
31'b0000000000000010000000000001010,
31'b1100010001010000000000000000000,
31'b0001000001010000000000000010010,
31'b0100000000100000000100100000000,
31'b0100000000100010000100100000000,
31'b0000110000100000100000000000000,
31'b0000010000010000000010001000000,
31'b0000000000010000000000000001010,
31'b0000000010100001000010000000000,
31'b1100010001100000000000000000000,
31'b0011001000000000000000001000100,
31'b0100000000010000000100100000000,
31'b0100000000100000000011000010000,
31'b0000110000010000100000000000000,
31'b0000100000000001000000000000110,
31'b0000000000100000000000000001010,
31'b0000000010010001000010000000000,
31'b0100000000000100000100100000000,
31'b0100010100000000000010000100000,
31'b0100000000000000000100100000000,
31'b0100000000000010000100100000000,
31'b0000110000000000100000000000000,
31'b0000110000000010100000000000000,
31'b0000000000000000001000001000100,
31'b0000000010000001000010000000000,
31'b1100010010000000000000000000000,
31'b0001000010000000000000000010010,
31'b1100010010000100000000000000000,
31'b0011000000000000000100000000101,
31'b1100010010001000000000000000000,
31'b0001000010001000000000000010010,
31'b1000000100000001000000000100000,
31'b1001000010000000000010000000001,
31'b1100010010010000000000000000000,
31'b0001000010010000000000000010010,
31'b1100000000100001000000001000000,
31'b0011000000001000000000000100010,
31'b0001001000000000000000100001010,
31'b0001000000000000000110010000000,
31'b1010000010100000010000000000000,
31'b0011000000000000000000000100010,
31'b1000000000000000010000000110000,
31'b1100100000000000001000000000010,
31'b1100000000010001000000001000000,
31'b0010000100001000000000000001001,
31'b1110000100000000000001000000000,
31'b0010000100000100000000000001001,
31'b1010000010010000010000000000000,
31'b0010000100000000000000000001001,
31'b1100000000000101000000001000000,
31'b0010000000001000100001010000000,
31'b1100000000000001000000001000000,
31'b0010000000000000000000101000100,
31'b1010000010000100010000000000000,
31'b0010000000000000100001010000000,
31'b1010000010000000010000000000000,
31'b0000000001000001000010000000000,
31'b1100010011000000000000000000000,
31'b0001000100000000100100001000000,
31'b0100001000000001000000010000000,
31'b0100001000000011000000010000000,
31'b0000010000000001001000000000100,
31'b0000010010000000000010001000000,
31'b0000000010000000000000000001010,
31'b0000000010000010000000000001010,
31'b0010100100000000100001000000000,
31'b0000000100000000010010000010000,
31'b0100001000010001000000010000000,
31'b0000001000000000000000100010010,
31'b0000100000000000000010000001100,
31'b0000000000000000101000000000010,
31'b0000000010010000000000000001010,
31'b0000000000100001000010000000000,
31'b1100000000000000000000110000001,
31'b0010000100000000000011001000000,
31'b0100001000100001000000010000000,
31'b0000000000011001000010000000000,
31'b0000110010010000100000000000000,
31'b0000000000010101000010000000000,
31'b0000000010100000000000000001010,
31'b0000000000010001000010000000000,
31'b0101010000000001000000000000001,
31'b0000000100000000100000100000001,
31'b0100000010000000000100100000000,
31'b0000000000001001000010000000000,
31'b0000110010000000100000000000000,
31'b0000000000000101000010000000000,
31'b0000000000000011000010000000000,
31'b0000000000000001000010000000000,
31'b1100010100000000000000000000000,
31'b0001000100000000000000000010010,
31'b1100010100000100000000000000000,
31'b0001001000100000100000000000001,
31'b1100010100001000000000000000000,
31'b0001000100001000000000000010010,
31'b1000000010000001000000000100000,
31'b1001000100000000000010000000001,
31'b1010000000000001000000000010000,
31'b0000010000000000100000010000000,
31'b1010000000000101000000000010000,
31'b0000101000000000000001000010000,
31'b1010000000001001000000000010000,
31'b0000010000001000100000010000000,
31'b1010000100100000010000000000000,
31'b0100100000000000000100110000000,
31'b1100010100100000000000000000000,
31'b0001001000000100100000000000001,
31'b0001001000000010100000000000001,
31'b0001001000000000100000000000001,
31'b1110000010000000000001000000000,
31'b0010000010000100000000000001001,
31'b1010000100010000010000000000000,
31'b0010000010000000000000000001001,
31'b1010000000100001000000000010000,
31'b0000010000100000100000010000000,
31'b1100000000000000000001000110000,
31'b0001010000000000000001000100010,
31'b1000010000000000000000001100000,
31'b1010000000000000000100010001000,
31'b1010000100000000010000000000000,
31'b1010000100000010010000000000000,
31'b1100010101000000000000000000000,
31'b0001000101000000000000000010010,
31'b0100000000000000001000000100100,
31'b0100000100000000000011000010000,
31'b0000011000000000000000010100000,
31'b0000010100000000000010001000000,
31'b0000000100000000000000000001010,
31'b0010000000000000010010000100000,
31'b1010000001000001000000000010000,
31'b0000010001000000100000010000000,
31'b0100000100100000000100100000000,
31'b1010100000000000010000010000000,
31'b0001101000000000000001000001000,
31'b0000010100010000000010001000000,
31'b0001000000100000000000000100001,
31'b1011000000000001000000000001000,
31'b0011000010000000000000000010001,
31'b1100000000000000001001100000000,
31'b0001000000000000000100000000110,
31'b1000101000000000001000000000100,
31'b0001100000000000000000010010010,
31'b1100110000000000000000010000000,
31'b0001000000010000000000000100001,
31'b0010000011000000000000000001001,
31'b0100010000000010000010000100000,
31'b0100010000000000000010000100000,
31'b0100000100000000000100100000000,
31'b0100010000000100000010000100000,
31'b0001000000000100000000000100001,
31'b0101100000000001000000100000000,
31'b0001000000000000000000000100001,
31'b0001000000000010000000000100001,
31'b1100010110000000000000000000000,
31'b0001000110000000000000000010010,
31'b1000000000001001000000000100000,
31'b1000010000000000100100000000001,
31'b1000000000000101000000000100000,
31'b1100100000000000000000100000001,
31'b1000000000000001000000000100000,
31'b1000000000000011000000000100000,
31'b1010000010000001000000000010000,
31'b0000010010000000100000010000000,
31'b1000010000000000010001000000000,
31'b1000010000000010010001000000000,
31'b1100000000000000010000001010000,
31'b0001010000000000010000001000010,
31'b1000000000010001000000000100000,
31'b1000000001000000010000000000011,
31'b1110000000001000000001000000000,
31'b0010000001000000000011001000000,
31'b1010010000000000000000001010000,
31'b0010000000001000000000000001001,
31'b1110000000000000000001000000000,
31'b0010000000000100000000000001001,
31'b1000000000100001000000000100000,
31'b0010000000000000000000000001001,
31'b0001100001000000000110000000000,
31'b0000000001000000100000100000001,
31'b1100000100000001000000001000000,
31'b0010000100000000000000101000100,
31'b1110000000010000000001000000000,
31'b0010000100000000100001010000000,
31'b1010000110000000010000000000000,
31'b0010000000010000000000000001001,
31'b0011000000100000000000000010001,
31'b0001000000000000100100001000000,
31'b1000011000000000000000000000110,
31'b1000001000010001100000000000000,
31'b1100000000000000001000010000010,
31'b0001010000000000001000010010000,
31'b1000000001000001000000000100000,
31'b1000000001000011000000000100000,
31'b0010100000000000100001000000000,
31'b0000000000000000010010000010000,
31'b1000010001000000010001000000000,
31'b1000001000000001100000000000000,
31'b0110000000000000001000000010100,
31'b0000000100000000101000000000010,
31'b1000000001010001000000000100000,
31'b1000000000000000010000000000011,
31'b0011000000000000000000000010001,
31'b0010000000000000000011001000000,
31'b0011000000000100000000000010001,
31'b0010000001001000000000000001001,
31'b1110000001000000000001000000000,
31'b0010000001000100000000000001001,
31'b1011000000000000000010000000010,
31'b0010000001000000000000000001001,
31'b0001100000000000000110000000000,
31'b0000000000000000100000100000001,
31'b0100100000000001100000000100000,
31'b0000000100001001000010000000000,
31'b0001100000001000000110000000000,
31'b0000000100000101000010000000000,
31'b0001000010000000000000000100001,
31'b0000000100000001000010000000000,
31'b1100011000000000000000000000000,
31'b0001001000000000000000000010010,
31'b1100011000000100000000000000000,
31'b0001001000000100000000000010010,
31'b1100011000001000000000000000000,
31'b0010100000000001000000001010000,
31'b1000000000000000001000010000100,
31'b1001001000000000000010000000001,
31'b1100011000010000000000000000000,
31'b0001001000010000000000000010010,
31'b0010000100000000110010000000000,
31'b0000100100000000000001000010000,
31'b0010000000000100001000000010010,
31'b1100000000000000010000000000101,
31'b0010000000000000001000000010010,
31'b0110100000000000010000000100000,
31'b0101000010000000000100000000000,
31'b0000110000000000000000000100000,
31'b0101000010000100000100000000000,
31'b0001000100000000100000000000001,
31'b0101000010001000000100000000000,
31'b0001000000000001000010100000000,
31'b1010001000010000010000000000000,
31'b0100100110000001000000000000000,
31'b0101000010010000000100000000000,
31'b0001000000000000000001010001000,
31'b1101000000000000000000010000001,
31'b0001000100010000100000000000001,
31'b1010001000000100010000000000000,
31'b1000010000000000000010010000000,
31'b1010001000000000010000000000000,
31'b1010001000000010010000000000000,
31'b1100011001000000000000000000000,
31'b0011000000100000000000001000100,
31'b0100000010000001000000010000000,
31'b0100001000000000000011000010000,
31'b0000010100000000000000010100000,
31'b0010000000000000000000100100010,
31'b0000001000000000000000000001010,
31'b0000001000000010000000000001010,
31'b1100000000000001000100000000001,
31'b0011000000000000001000000001010,
31'b0100001000100000000100100000000,
31'b0000000010000000000000100010010,
31'b0001100100000000000001000001000,
31'b1100010000000000100000000100000,
31'b0000001000010000000000000001010,
31'b0000001010100001000010000000000,
31'b0101000011000000000100000000000,
31'b0011000000000000000000001000100,
31'b0100001000010000000100100000000,
31'b1010000000000000110000000100000,
31'b0000111000010000100000000000000,
31'b0011000000001000000000001000100,
31'b0000001000100000000000000001010,
31'b0100000010000000000100000011000,
31'b0100010000000000000000011000000,
31'b0110000000000000000100000101000,
31'b0100001000000000000100100000000,
31'b0100001000000010000100100000000,
31'b0000111000000000100000000000000,
31'b1000010001000000000010010000000,
31'b0000000000000000000001010010000,
31'b0000001010000001000010000000000,
31'b0000000000000000001000000100010,
31'b0100100000000000010000000010000,
31'b0100000001000001000000010000000,
31'b0100100000000100010000000010000,
31'b0100000100000000000000000001100,
31'b0100100000001000010000000010000,
31'b1000001100000001000000000100000,
31'b1000000100000000000001000000101,
31'b0100000000000000000000101000001,
31'b0100100000010000010000000010000,
31'b0100000001010001000000010000000,
31'b0000100000000001000000001100000,
31'b0001000000000000000000100001010,
31'b1000000001000000000010100000001,
31'b0011010000000000010100000000000,
31'b0011001000000000000000000100010,
31'b0101000000000000000100000000000,
31'b0101000000000010000100000000000,
31'b0101000000000100000100000000000,
31'b0101000000000110000100000000000,
31'b0101000000001000000100000000000,
31'b0101000000001010000100000000000,
31'b0101000000001100000100000000000,
31'b0100100100000001000000000000000,
31'b0101000000010000000100000000000,
31'b0110100000000000000001001000000,
31'b1100001000000001000000001000000,
31'b0010110000001000000000000010000,
31'b0101000000011000000100000000000,
31'b1000010010000000000010010000000,
31'b1010001010000000010000000000000,
31'b0010110000000000000000000010000,
31'b0100000000000101000000010000000,
31'b0100100001000000010000000010000,
31'b0100000000000001000000010000000,
31'b0100000000000011000000010000000,
31'b0100000101000000000000000001100,
31'b1010000000000000100001001000000,
31'b0100000000001001000000010000000,
31'b0100000000100000000100000011000,
31'b0100000001000000000000101000001,
31'b0000000000000100000000100010010,
31'b0100000000010001000000010000000,
31'b0000000000000000000000100010010,
31'b1001100000000000100100000000000,
31'b1000000000000000000010100000001,
31'b0100000000011001000000010000000,
31'b0000001000100001000010000000000,
31'b0101000001000000000100000000000,
31'b0101000001000010000100000000000,
31'b0100000000100001000000010000000,
31'b0100000000100011000000010000000,
31'b1011000000000000010000100000000,
31'b1001000000000000000110001000000,
31'b0100000000101001000000010000000,
31'b0100000000000000000100000011000,
31'b0101000001010000000100000000000,
31'b1000000100000000001010000000010,
31'b0100001010000000000100100000000,
31'b0000001000001001000010000000000,
31'b1010100000000000000011000000000,
31'b1000000000000000110000000010000,
31'b0000001000000011000010000000000,
31'b0000001000000001000010000000000,
31'b1100011100000000000000000000000,
31'b0001001100000000000000000010010,
31'b0011000000000000000100001010000,
31'b0001000000100000100000000000001,
31'b0100000010000000000000000001100,
31'b0100110000010000000000001000000,
31'b1000001010000001000000000100000,
31'b1001000000000001001000000010000,
31'b1010001000000001000000000010000,
31'b0000100000000100000001000010000,
31'b0010000000000000110010000000000,
31'b0000100000000000000001000010000,
31'b0100110000000010000000001000000,
31'b0100110000000000000000001000000,
31'b0100100000000000000010000001010,
31'b0100000000000000101000000000100,
31'b0101000110000000000100000000000,
31'b0001000000000100100000000000001,
31'b0001000000000010100000000000001,
31'b0001000000000000100000000000001,
31'b0100010000000000100010000000000,
31'b0100100010000101000000000000000,
31'b0100100010000011000000000000000,
31'b0100100010000001000000000000000,
31'b0010000000000100000000100010001,
31'b0001000100000000000001010001000,
31'b0010000000000000000000100010001,
31'b0001000000010000100000000000001,
31'b1010000000000000000010100000010,
31'b1000010100000000000010010000000,
31'b1010001100000000010000000000000,
31'b0100100010010001000000000000000,
31'b1000000000000001001000000001000,
31'b1000010000100000100000001000000,
31'b1000010010000000000000000000110,
31'b1000100000100000001000000000100,
31'b0000010000000000000000010100000,
31'b0010000000000000000100001001000,
31'b0000010000000100000000010100000,
31'b0010001000000000010010000100000,
31'b1000110000000000000010000000000,
31'b1000110000000010000010000000000,
31'b1000110000000100000010000000000,
31'b1000000010000001100000000000000,
31'b0001100000000000000001000001000,
31'b0111000000000000000000000100100,
31'b0001100000000100000001000001000,
31'b1101100000000000000000000000001,
31'b1000010000000010100000001000000,
31'b1000010000000000100000001000000,
31'b1000100000000010001000000000100,
31'b1000100000000000001000000000100,
31'b0000010000100000000000010100000,
31'b1000010000001000100000001000000,
31'b0001010000000000100001000000010,
31'b1100000000000000100001000010000,
31'b1000110000100000000010000000000,
31'b1000010000010000100000001000000,
31'b0110000000000000010000010100000,
31'b1000100000010000001000000000100,
31'b0001100000100000000001000001000,
31'b0011000000000000000000100001001,
31'b0001001000000000000000000100001,
31'b0001000000000001000001000000100,
31'b0100000000001000000000000001100,
31'b0100100100000000010000000010000,
31'b1000010001000000000000000000110,
31'b1000000001010001100000000000000,
31'b0100000000000000000000000001100,
31'b0100000000000010000000000001100,
31'b1000001000000001000000000100000,
31'b1000000000000000000001000000101,
31'b0100000100000000000000101000001,
31'b1010000000000000000011010000000,
31'b1000011000000000010001000000000,
31'b1000000001000001100000000000000,
31'b0100000000010000000000000001100,
31'b0100110010000000000000001000000,
31'b1000001000010001000000000100000,
31'b1000000001001001100000000000000,
31'b0101000100000000000100000000000,
31'b0101000100000010000100000000000,
31'b0101000100000100000100000000000,
31'b0100100000001001000000000000000,
31'b0000000000000000000000100100001,
31'b0100100000000101000000000000000,
31'b0100100000000011000000000000000,
31'b0100100000000001000000000000000,
31'b0001000000000000001000000001001,
31'b1001000000000000100100010000000,
31'b0010010000000000010000000001100,
31'b1101000000000000001001000000000,
31'b0100000000000000001000001000010,
31'b0100100000010101000000000000000,
31'b0100100000010011000000000000000,
31'b0100100000010001000000000000000,
31'b1000010000000100000000000000110,
31'b1000000000010101100000000000000,
31'b1000010000000000000000000000110,
31'b1000000000010001100000000000000,
31'b0100000001000000000000000001100,
31'b0101100000000000000100010000000,
31'b1000010000001000000000000000110,
31'b1000000001000000000001000000101,
31'b1000110010000000000010000000000,
31'b1000000000000101100000000000000,
31'b1000000000000011100000000000000,
31'b1000000000000001100000000000000,
31'b0110000000000000000001011000000,
31'b1000000100000000000010100000001,
31'b1000010000000000000100000100001,
31'b1000000000001001100000000000000,
31'b0101000101000000000100000000000,
31'b1000010010000000100000001000000,
31'b1000100000000001000010001000000,
31'b1000100010000000001000000000100,
31'b0100000000000000010000010010000,
31'b0100100001000101000000000000000,
31'b0100100001000011000000000000000,
31'b0100100001000001000000000000000,
31'b1000100000000000100000000001100,
31'b1000000000000000001010000000010,
31'b1000010000000000001000001001000,
31'b1000000000100001100000000000000,
31'b0100000001000000001000001000010,
31'b0000000000000100001000000010001,
31'b0000000000000010001000000010001,
31'b0000000000000000001000000010001,
31'b1100100000000000000000000000000,
31'b0000001000100000000000000100000,
31'b1100100000000100000000000000000,
31'b0000100000000000000001000001001,
31'b1100100000001000000000000000000,
31'b0000100001000000000010001000000,
31'b1100100000001100000000000000000,
31'b0000100001000100000010001000000,
31'b1100100000010000000000000000000,
31'b0000100100000000100000010000000,
31'b1100100000010100000000000000000,
31'b0001010000000000000000010100001,
31'b0000000001100000100000000000000,
31'b0100001100000000000000001000000,
31'b0110000000000000000100000000010,
31'b0110000000000010000100000000010,
31'b0000001000000010000000000100000,
31'b0000001000000000000000000100000,
31'b0010000000000000000000100001000,
31'b0000001000000100000000000100000,
31'b0000000001010000100000000000000,
31'b0000001000001000000000000100000,
31'b0010000000001000000000100001000,
31'b0000001000001100000000000100000,
31'b0000000001001000100000000000000,
31'b0000001000010000000000000100000,
31'b0010000000010000000000100001000,
31'b0001000000000000100000000011000,
31'b0000000001000000100000000000000,
31'b0000000001000010100000000000000,
31'b0000000001000100100000000000000,
31'b0010001010000000000000000010000,
31'b1100100001000000000000000000000,
31'b0000100000001000000010001000000,
31'b1100100001000100000000000000000,
31'b0000100001000000000001000001001,
31'b0000000000110000100000000000000,
31'b0000100000000000000010001000000,
31'b0000110000000000000000000001010,
31'b0000100000000100000010001000000,
31'b0000000000101000100000000000000,
31'b1000000000000000000000011100000,
31'b1000000000000000010000100000010,
31'b1000000000000100000000011100000,
31'b0000000000100000100000000000000,
31'b0000000000100010100000000000000,
31'b0000000000100100100000000000000,
31'b0000000010000000000000001000110,
31'b0000000000011000100000000000000,
31'b0000001001000000000000000100000,
31'b0010000001000000000000100001000,
31'b0000001001000100000000000100000,
31'b0000000000010000100000000000000,
31'b0000000000010010100000000000000,
31'b0000000000010100100000000000000,
31'b0000000010000000001000000001000,
31'b0000000000001000100000000000000,
31'b0000000000001010100000000000000,
31'b0000000000001100100000000000000,
31'b0001000010000000000000100100000,
31'b0000000000000000100000000000000,
31'b0000000000000010100000000000000,
31'b0000000000000100100000000000000,
31'b0000000000000110100000000000000,
31'b1100100010000000000000000000000,
31'b0000100000000000011100000000000,
31'b1100100010000100000000000000000,
31'b0000100010000000000001000001001,
31'b1100100010001000000000000000000,
31'b0000100011000000000010001000000,
31'b0001001000100000100000100000000,
31'b0000001000000000010001001000000,
31'b1100100010010000000000000000000,
31'b0010001100000001010000000000000,
31'b1100000000000000000010000000110,
31'b0010001000101000000000000010000,
31'b0100000000000000000000000010101,
31'b0100001110000000000000001000000,
31'b0110000010000000000100000000010,
31'b0010001000100000000000000010000,
31'b0001000000000000001000000010000,
31'b0000001010000000000000000100000,
31'b0010000010000000000000100001000,
31'b0000001010000100000000000100000,
31'b0001000000001000001000000010000,
31'b0000001010001000000000000100000,
31'b0001001000000000100000100000000,
31'b0000000001000000001000000001000,
31'b0001000000010000001000000010000,
31'b0010000000000000101000100000000,
31'b0010001000001010000000000010000,
31'b0010001000001000000000000010000,
31'b0000000011000000100000000000000,
31'b0010001000000100000000000010000,
31'b0010001000000010000000000010000,
31'b0010001000000000000000000010000,
31'b1100100011000000000000000000000,
31'b0000100010001000000010001000000,
31'b0010010000000000000000010001001,
31'b0000000000101000001000000001000,
31'b0000100000000001001000000000100,
31'b0000100010000000000010001000000,
31'b0000010000000001100000001000000,
31'b0000000000100000001000000001000,
31'b1001000000000000000001000000100,
31'b1001000000000010000001000000100,
31'b1001000000000100000001000000100,
31'b0001000000100000000000100100000,
31'b0000000010100000100000000000000,
31'b0000000010100010100000000000000,
31'b0000000010100100100000000000000,
31'b0000000000000000000000001000110,
31'b0001000001000000001000000010000,
31'b0000001011000000000000000100000,
31'b0010000000000000100000000110000,
31'b0000000000001000001000000001000,
31'b0000000010010000100000000000000,
31'b0000000000000100001000000001000,
31'b0000000000000010001000000001000,
31'b0000000000000000001000000001000,
31'b0000000010001000100000000000000,
31'b0001000000000100000000100100000,
31'b0001000000000010000000100100000,
31'b0001000000000000000000100100000,
31'b0000000010000000100000000000000,
31'b0000000010000010100000000000000,
31'b0000000010000100100000000000000,
31'b0000000000010000001000000001000,
31'b1100100100000000000000000000000,
31'b0000100000010000100000010000000,
31'b1100100100000100000000000000000,
31'b0000100100000000000001000001001,
31'b1100100100001000000000000000000,
31'b1000000000000000100010000100000,
31'b0011000000000000000100100000100,
31'b1101000000000001000100000000000,
31'b1000001001000000000010000000000,
31'b0000100000000000100000010000000,
31'b1000100010000000010001000000000,
31'b0000100000000100100000010000000,
31'b0100001000000010000000001000000,
31'b0100001000000000000000001000000,
31'b0110000100000000000100000000010,
31'b0100001000000100000000001000000,
31'b0000000000000000000010011000000,
31'b0000001100000000000000000100000,
31'b0010000100000000000000100001000,
31'b0000010000000000000000010001010,
31'b0000000101010000100000000000000,
31'b1100000001000000000000010000000,
31'b0010000100001000000000100001000,
31'b1100000001000100000000010000000,
31'b0000000101001000100000000000000,
31'b0000100000100000100000010000000,
31'b0010000100010000000000100001000,
31'b0001100000000000000001000100010,
31'b0000000101000000100000000000000,
31'b0100001000100000000000001000000,
31'b0010000000000000000000001000101,
31'b0100001000100100000000001000000,
31'b1000001000010000000010000000000,
31'b1100000000101000000000010000000,
31'b1101000000000000010000000000100,
31'b0011000000000001010000100000000,
31'b0000101000000000000000010100000,
31'b1100000000100000000000010000000,
31'b0000110100000000000000000001010,
31'b1100000000100100000000010000000,
31'b1000001000000000000010000000000,
31'b1000001000000010000010000000000,
31'b1000001000000100000010000000000,
31'b1010010000000000010000010000000,
31'b0000000100100000100000000000000,
31'b0100001001000000000000001000000,
31'b0000001000000000000000000010011,
31'b0100001001000100000000001000000,
31'b0000000100011000100000000000000,
31'b1100000000001000000000010000000,
31'b0010000101000000000000100001000,
31'b1100000000001100000000010000000,
31'b0000000100010000100000000000000,
31'b1100000000000000000000010000000,
31'b0000000100010100100000000000000,
31'b1100000000000100000000010000000,
31'b0000000100001000100000000000000,
31'b0100100000000000000010000100000,
31'b0000000100001100100000000000000,
31'b0100100000000100000010000100000,
31'b0000000100000000100000000000000,
31'b0000000100000010100000000000000,
31'b0000000100000100100000000000000,
31'b0100000010000000000100000000001,
31'b1100100110000000000000000000000,
31'b0010001000010001010000000000000,
31'b1001000000000000000010100000000,
31'b1001000000000010000010100000000,
31'b0010010000000001000000000000101,
31'b1100010000000000000000100000001,
31'b0001000000000001011000000000000,
31'b0101000001000000000000101000000,
31'b1000100000000100010001000000000,
31'b0010001000000001010000000000000,
31'b1000100000000000010001000000000,
31'b1010000000000000100010000010000,
31'b0100001010000010000000001000000,
31'b0100001010000000000000001000000,
31'b1000100000001000010001000000000,
31'b0100001010000100000000001000000,
31'b0001000100000000001000000010000,
31'b0000001110000000000000000100000,
31'b1010100000000000000000001010000,
31'b0100011000001001000000000000000,
31'b0001000100001000001000000010000,
31'b1100000011000000000000010000000,
31'b0100011000000011000000000000000,
31'b0100011000000001000000000000000,
31'b0001010001000000000110000000000,
31'b0010001000100001010000000000000,
31'b1000100000100000010001000000000,
31'b1010000000000000010000100000001,
31'b0000000111000000100000000000000,
31'b0100001010100000000000001000000,
31'b0100001000000000100000000000110,
31'b0100000001000000000100000000001,
31'b1100000000000000000001100000010,
31'b0010010000000000010100000000001,
31'b1001000001000000000010100000000,
31'b0001000000000000001100000000100,
31'b0010001000010000000100000000100,
31'b1100000010100000000000010000000,
31'b0101000000000010000000101000000,
31'b0101000000000000000000101000000,
31'b1000001010000000000010000000000,
31'b1000001010000010000010000000000,
31'b1000100001000000010001000000000,
31'b0100000000101000000100000000001,
31'b0010001000000000000100000000100,
31'b0100001011000000000000001000000,
31'b0110000000000000100000001010000,
31'b0100000000100000000100000000001,
31'b0001010000010000000110000000000,
31'b1100000010001000000000010000000,
31'b0100000000001000110001000000000,
31'b0100000000000000000000000100110,
31'b0000000110010000100000000000000,
31'b1100000010000000000000010000000,
31'b0100000000000000110001000000000,
31'b0000000100000000001000000001000,
31'b0001010000000000000110000000000,
31'b0100100010000000000010000100000,
31'b0100010000000001100000000100000,
31'b0100000000001000000100000000001,
31'b0000000110000000100000000000000,
31'b0100000000000100000100000000001,
31'b0100000000000010000100000000001,
31'b0100000000000000000100000000001,
31'b0000000000100010000000000100000,
31'b0000000000100000000000000100000,
31'b1000000000000000000001100000100,
31'b0000000000100100000000000100000,
31'b1000000000000000100000011000000,
31'b0000000000101000000000000100000,
31'b1000000000001000000001100000100,
31'b0000000010000000010001001000000,
31'b1000000101000000000010000000000,
31'b0000000000110000000000000100000,
31'b1000000101000100000010000000000,
31'b0000010100000000000001000010000,
31'b0100000100000010000000001000000,
31'b0100000100000000000000001000000,
31'b0110001000000000000100000000010,
31'b0100000100000100000000001000000,
31'b0000000000000010000000000100000,
31'b0000000000000000000000000100000,
31'b0000000000000110000000000100000,
31'b0000000000000100000000000100000,
31'b0000000000001010000000000100000,
31'b0000000000001000000000000100000,
31'b0001000010000000100000100000000,
31'b0000000000001100000000000100000,
31'b0000000000010010000000000100000,
31'b0000000000010000000000000100000,
31'b0000000001000000001000100010000,
31'b0000000000010100000000000100000,
31'b0000001001000000100000000000000,
31'b0000000000011000000000000100000,
31'b0010000010000010000000000010000,
31'b0010000010000000000000000010000,
31'b1000000100010000000010000000000,
31'b0000000001100000000000000100000,
31'b1000000100010100000010000000000,
31'b0000000001100100000000000100000,
31'b0000100100000000000000010100000,
31'b0000101000000000000010001000000,
31'b0001010000000000100000010000001,
31'b0000101000000100000010001000000,
31'b1000000100000000000010000000000,
31'b1000000100000010000010000000000,
31'b1000000100000100000010000000000,
31'b1000010000000000000100100100000,
31'b0000001000100000100000000000000,
31'b0100000101000000000000001000000,
31'b0000001000100100100000000000000,
31'b0110000000000000100000000000101,
31'b0000000001000010000000000100000,
31'b0000000001000000000000000100000,
31'b0000000001000110000000000100000,
31'b0000000001000100000000000100000,
31'b0000001000010000100000000000000,
31'b0000000001001000000000000100000,
31'b0001000000000000000000000111000,
31'b0000001010000000001000000001000,
31'b0000001000001000100000000000000,
31'b0000000001010000000000000100000,
31'b0000000000000000001000100010000,
31'b0000000001010100000000000100000,
31'b0000001000000000100000000000000,
31'b0000001000000010100000000000000,
31'b0000001000000100100000000000000,
31'b0010000011000000000000000010000,
31'b1001000000000000010000000000010,
31'b0000000010100000000000000100000,
31'b1001000000000100010000000000010,
31'b0000000010100100000000000100000,
31'b1001000000001000010000000000010,
31'b0000000010101000000000000100000,
31'b0001000000100000100000100000000,
31'b0000000000000000010001001000000,
31'b1001000000010000010000000000010,
31'b0010000100000001010000000000000,
31'b0010000000101010000000000010000,
31'b0010000000101000000000000010000,
31'b0100001000000000000000000010101,
31'b0100000110000000000000001000000,
31'b0010000000100010000000000010000,
31'b0010000000100000000000000010000,
31'b0000000010000010000000000100000,
31'b0000000010000000000000000100000,
31'b0001000000001000100000100000000,
31'b0000000010000100000000000100000,
31'b0001000000000100100000100000000,
31'b0000000010001000000000000100000,
31'b0001000000000000100000100000000,
31'b0010000000010000000000000010000,
31'b0011000001000000000000000001000,
31'b0000000010010000000000000100000,
31'b0010000000001010000000000010000,
31'b0010000000001000000000000010000,
31'b0010000000000110000000000010000,
31'b0010000000000100000000000010000,
31'b0010000000000010000000000010000,
31'b0010000000000000000000000010000,
31'b1001000001000000010000000000010,
31'b0000000011100000000000000100000,
31'b1100000000000000010011000000000,
31'b0000001000101000001000000001000,
31'b0010000100010000000100000000100,
31'b0000101010000000000010001000000,
31'b0101010000000000010000000001000,
31'b0000001000100000001000000001000,
31'b1000000110000000000010000000000,
31'b1001000000000001000000000100001,
31'b1101100000000000000000100000000,
31'b0011100000000001000000000000100,
31'b0010000100000000000100000000100,
31'b0100000111000000000000001000000,
31'b0010000100000100000100000000100,
31'b0010000001100000000000000010000,
31'b0011000000010000000000000001000,
31'b0000000011000000000000000100000,
31'b0011000000010100000000000001000,
31'b0000001000001000001000000001000,
31'b0010000000000000001000100100000,
31'b0000001000000100001000000001000,
31'b0001000001000000100000100000000,
31'b0000001000000000001000000001000,
31'b0011000000000000000000000001000,
31'b0011000000000010000000000001000,
31'b0011000000000100000000000001000,
31'b0010000001001000000000000010000,
31'b0000001010000000100000000000000,
31'b0010000001000100000000000010000,
31'b0010000001000010000000000010000,
31'b0010000001000000000000000010000,
31'b1000000001010000000010000000000,
31'b0000000100100000000000000100000,
31'b1000000100000000000001100000100,
31'b0000010000010000000001000010000,
31'b0100000000010010000000001000000,
31'b0100000000010000000000001000000,
31'b0100100000000001001000000000010,
31'b0100000000010100000000001000000,
31'b1000000001000000000010000000000,
31'b0100000000001000000000001000000,
31'b1000000001000100000010000000000,
31'b0000010000000000000001000010000,
31'b0100000000000010000000001000000,
31'b0100000000000000000000001000000,
31'b0100000000000110000000001000000,
31'b0100000000000100000000001000000,
31'b0000000100000010000000000100000,
31'b0000000100000000000000000100000,
31'b0000010000000000000110100000000,
31'b0000000100000100000000000100000,
31'b0100100000000000100010000000000,
31'b0000000100001000000000000100000,
31'b0100100000000100100010000000000,
31'b0100010010000001000000000000000,
31'b1000000001100000000010000000000,
31'b0000000100010000000000000100000,
31'b1000000001100100000010000000000,
31'b0000010000100000000001000010000,
31'b0100000000100010000000001000000,
31'b0100000000100000000000001000000,
31'b0100000010000000100000000000110,
31'b0100000000100100000000001000000,
31'b1000000000010000000010000000000,
31'b1000000000010010000010000000000,
31'b1000000000010100000010000000000,
31'b1000010000100000001000000000100,
31'b0000100000000000000000010100000,
31'b0100000001010000000000001000000,
31'b0000100000000100000000010100000,
31'b0100000001010100000000001000000,
31'b1000000000000000000010000000000,
31'b1000000000000010000010000000000,
31'b1000000000000100000010000000000,
31'b1000000000000110000010000000000,
31'b1000000000001000000010000000000,
31'b0100000001000000000000001000000,
31'b0000000000000000000000000010011,
31'b0100000001000100000000001000000,
31'b1000000000110000000010000000000,
31'b0000000101000000000000000100000,
31'b1000010000000010001000000000100,
31'b1000010000000000001000000000100,
31'b0000100000100000000000010100000,
31'b1100001000000000000000010000000,
31'b0001100000000000100001000000010,
31'b1100001000000100000000010000000,
31'b1000000000100000000010000000000,
31'b1000000000100010000010000000000,
31'b1000000000100100000010000000000,
31'b1000010000010000001000000000100,
31'b0000001100000000100000000000000,
31'b0100000001100000000000001000000,
31'b0000001100000100100000000000000,
31'b0100001010000000000100000000001,
31'b1001000100000000010000000000010,
31'b0010000000010001010000000000000,
31'b1001001000000000000010100000000,
31'b0110000000000000000000001110000,
31'b0100110000000000000000000001100,
31'b0100000010010000000000001000000,
31'b0100010000100011000000000000000,
31'b0100010000100001000000000000000,
31'b1000000011000000000010000000000,
31'b0010000000000001010000000000000,
31'b1000101000000000010001000000000,
31'b0010000000000101010000000000000,
31'b0100000010000010000000001000000,
31'b0100000010000000000000001000000,
31'b0100000010000110000000001000000,
31'b0100000010000100000000001000000,
31'b0001000000000001000010000000001,
31'b0000000110000000000000000100000,
31'b0100010000001011000000000000000,
31'b0100010000001001000000000000000,
31'b0100100010000000100010000000000,
31'b0100010000000101000000000000000,
31'b0100010000000011000000000000000,
31'b0100010000000001000000000000000,
31'b1000000011100000000010000000000,
31'b0010000000100001010000000000000,
31'b0100000000001000100000000000110,
31'b0100000000000000010001000100000,
31'b0100000010100010000000001000000,
31'b0100000010100000000000001000000,
31'b0100000000000000100000000000110,
31'b0010000100000000000000000010000,
31'b1000000010010000000010000000000,
31'b1000000010010010000010000000000,
31'b1000100000000000000000000000110,
31'b1000100000000010000000000000110,
31'b0010000000010000000100000000100,
31'b0101010000000000000100010000000,
31'b1010000000000000000010000110000,
31'b0101001000000000000000101000000,
31'b1000000010000000000010000000000,
31'b1000000010000010000010000000000,
31'b1000000010000100000010000000000,
31'b1000110000000001100000000000000,
31'b0010000000000000000100000000100,
31'b0100000011000000000000001000000,
31'b0010000000000100000100000000100,
31'b0100001000100000000100000000001,
31'b1000000010110000000010000000000,
31'b1000000000000001000000000001010,
31'b1000100000100000000000000000110,
31'b1000010010000000001000000000100,
31'b0010000100000000001000100100000,
31'b1100001010000000000000010000000,
31'b0100010001000011000000000000000,
31'b0100010001000001000000000000000,
31'b1000000010100000000010000000000,
31'b1000000010100010000010000000000,
31'b1000100000000000001000001001000,
31'b0100001000001000000100000000001,
31'b0010000000100000000100000000100,
31'b0100001000000100000100000000001,
31'b0100001000000010000100000000001,
31'b0100001000000000000100000000001,
31'b1100110000000000000000000000000,
31'b0001100000000000000000000010010,
31'b1100110000000100000000000000000,
31'b0001100000000100000000000010010,
31'b1100110000001000000000000000000,
31'b0011000000000000000010000100100,
31'b1000000000000000100100100000000,
31'b1001100000000000000010000000001,
31'b1100110000010000000000000000000,
31'b0001100000010000000000000010010,
31'b0001000000000010000000010100001,
31'b0001000000000000000000010100001,
31'b0100000000000000010000100001000,
31'b0100011100000000000000001000000,
31'b1010100000100000010000000000000,
31'b1011000000000000000100000010000,
31'b0000000000000000010100000000010,
31'b0000011000000000000000000100000,
31'b0010010000000000000000100001000,
31'b0000011000000100000000000100000,
31'b0000010001010000100000000000000,
31'b0000011000001000000000000100000,
31'b1010100000010000010000000000000,
31'b0100001110000001000000000000000,
31'b0000010001001000100000000000000,
31'b0000011000010000000000000100000,
31'b1100000000000000100000000001010,
31'b0001010000000000100000000011000,
31'b0000010001000000100000000000000,
31'b0000010001000010100000000000000,
31'b1010100000000000010000000000000,
31'b1010100000000010010000000000000,
31'b1100110001000000000000000000000,
31'b0001100001000000000000000010010,
31'b0110000000000000110000000000000,
31'b0110000000000010110000000000000,
31'b0000100000000100000000000001010,
31'b0000110000000000000010001000000,
31'b0000100000000000000000000001010,
31'b0000100000000010000000000001010,
31'b1010000000000000000100000001000,
31'b1010000000000010000100000001000,
31'b1010000000000100000100000001000,
31'b1010000100000000010000010000000,
31'b0000010000100000100000000000000,
31'b0000010000100010100000000000000,
31'b0000100000010000000000000001010,
31'b0000100010100001000010000000000,
31'b0000010000011000100000000000000,
31'b0000011001000000000000000100000,
31'b0110000000100000110000000000000,
31'b1000001100000000001000000000100,
31'b0000010000010000100000000000000,
31'b0000000000000001000000000000110,
31'b0000100000100000000000000001010,
31'b0000010010000000001000000001000,
31'b0000010000001000100000000000000,
31'b0000010000001010100000000000000,
31'b0100100000000000000100100000000,
31'b0101000000000000100010000000001,
31'b0000010000000000100000000000000,
31'b0000010000000010100000000000000,
31'b0000010000000100100000000000000,
31'b0000100010000001000010000000000,
31'b1100110010000000000000000000000,
31'b1001000000000000000100000100000,
31'b0010000001000000000000010001001,
31'b1100000000000001100010000000000,
31'b0010000100000001000000000000101,
31'b1100000100000000000000100000001,
31'b0000000100000000000001100001000,
31'b0100001100100001000000000000000,
31'b0010000101000000100001000000000,
31'b1100000000000000000000001001100,
31'b0000000100000001000010010000000,
31'b0001000000000000000010000010100,
31'b0000000001000000000010000001100,
31'b1001000000000000000000000000111,
31'b0000000100010000000001100001000,
31'b0011100000000000000000000100010,
31'b0001010000000000001000000010000,
31'b1100000000000000001000000000010,
31'b0010010010000000000000100001000,
31'b1100000000000100001000000000010,
31'b0001010000001000001000000010000,
31'b1100000000001000001000000000010,
31'b0101000000000000001001001000000,
31'b0100001100000001000000000000000,
31'b0001010000010000001000000010000,
31'b1100000000010000001000000000010,
31'b1100100000000001000000001000000,
31'b0010100000000000000000101000100,
31'b0000010011000000100000000000000,
31'b0010100000000000100001010000000,
31'b1010100010000000010000000000000,
31'b0010011000000000000000000010000,
31'b0010000100010000100001000000000,
31'b1110000000000000000001010000000,
31'b0010000000000000000000010001001,
31'b1010000000000000101100000000000,
31'b0000000000010000000010000001100,
31'b0000110010000000000010001000000,
31'b0000000000000001100000001000000,
31'b0000010000100000001000000001000,
31'b0010000100000000100001000000000,
31'b0110000000000000011000000001000,
31'b0010000100000100100001000000000,
31'b0001010000100000000000100100000,
31'b0000000000000000000010000001100,
31'b0000100000000000101000000000010,
31'b0000000000010001100000001000000,
31'b0000100000100001000010000000000,
31'b0001010001000000001000000010000,
31'b1100000001000000001000000000010,
31'b1000000000000011000000010100000,
31'b1000000000000001000000010100000,
31'b0000010010010000100000000000000,
31'b0000010000000100001000000001000,
31'b0000010000000010001000000001000,
31'b0000010000000000001000000001000,
31'b0001000100000000000110000000000,
31'b0001010000000100000000100100000,
31'b0100100010000000000100100000000,
31'b0001010000000000000000100100000,
31'b0000010010000000100000000000000,
31'b0000100000000101000010000000000,
31'b0000100000000011000010000000000,
31'b0000100000000001000010000000000,
31'b1100110100000000000000000000000,
31'b0001100100000000000000000010010,
31'b0000001000100000000110100000000,
31'b0000001000010000000001000010000,
31'b0011000000000000001001000010000,
31'b1100000010000000000000100000001,
31'b0000000010000000000001100001000,
31'b0100001010100001000000000000000,
31'b1010100000000001000000000010000,
31'b0000110000000000100000010000000,
31'b0000001000000010000001000010000,
31'b0000001000000000000001000010000,
31'b0100011000000010000000001000000,
31'b0100011000000000000000001000000,
31'b0100001000000000000010000001010,
31'b0100000000000000000100110000000,
31'b0000010000000000000010011000000,
31'b0000011100000000000000000100000,
31'b0000001000000000000110100000000,
31'b0000000000000000000000010001010,
31'b0001000001000000000000010010010,
31'b1100010001000000000000010000000,
31'b0100001010000011000000000000000,
31'b0100001010000001000000000000000,
31'b0001000011000000000110000000000,
31'b0000110000100000100000010000000,
31'b0100000010000000000101000000010,
31'b0000001000100000000001000010000,
31'b0001000000000000011000001000000,
31'b0101000001000001000000100000000,
31'b1010100100000000010000000000000,
31'b0100001010010001000000000000000,
31'b1110000000000000001000000000001,
31'b0010000010000000010100000000001,
31'b0110000100000000110000000000000,
31'b0010000000000000001001000001000,
31'b0001001000010000000001000001000,
31'b1100010000100000000000010000000,
31'b0000100100000000000000000001010,
31'b0010100000000000010010000100000,
31'b1000011000000000000010000000000,
31'b1010000000000100010000010000000,
31'b1010000000000010010000010000000,
31'b1010000000000000010000010000000,
31'b0001001000000000000001000001000,
31'b0101000000100001000000100000000,
31'b0001100000100000000000000100001,
31'b1101001000000000000000000000001,
31'b0001000010010000000110000000000,
31'b1100010000001000000000010000000,
31'b1001000000000000000010010000001,
31'b1000001000000000001000000000100,
31'b0001000000000000000000010010010,
31'b1100010000000000000000010000000,
31'b0001100000010000000000000100001,
31'b1100010000000100000000010000000,
31'b0001000010000000000110000000000,
31'b0101000000001001000000100000000,
31'b0100100100000000000100100000000,
31'b1010000000100000010000010000000,
31'b0000010100000000100000000000000,
31'b0101000000000001000000100000000,
31'b0001100000000000000000000100001,
31'b0101000000000101000000100000000,
31'b0010000001010000100001000000000,
31'b1100000000001000000000100000001,
31'b0000000000010001000010010000000,
31'b0100001000101001000000000000000,
31'b0010000000000001000000000000101,
31'b1100000000000000000000100000001,
31'b0000000000000000000001100001000,
31'b0100001000100001000000000000000,
31'b0010000001000000100001000000000,
31'b0010011000000001010000000000000,
31'b0000000000000001000010010000000,
31'b0000001010000000000001000010000,
31'b0010000001001000100001000000000,
31'b1100000000010000000000100000001,
31'b0000000000010000000001100001000,
31'b0100001000110001000000000000000,
31'b0001010100000000001000000010000,
31'b1100000100000000001000000000010,
31'b0100001000001011000000000000000,
31'b0100001000001001000000000000000,
31'b1110100000000000000001000000000,
31'b1000000000000000000000000101100,
31'b0100001000000011000000000000000,
31'b0100001000000001000000000000000,
31'b0001000001000000000110000000000,
31'b1001000000000000001000100000100,
31'b0100000000000000000101000000010,
31'b0100001000011001000000000000000,
31'b0001000010000000011000001000000,
31'b1101000000000000000100001000000,
31'b0100001000010011000000000000000,
31'b0100001000010001000000000000000,
31'b0010000000010000100001000000000,
31'b0010000000000000010100000000001,
31'b0010000100000000000000010001001,
31'b0010000010000000001001000001000,
31'b0010000001000001000000000000101,
31'b1100000001000000000000100000001,
31'b0000000100000001100000001000000,
31'b0101010000000000000000101000000,
31'b0010000000000000100001000000000,
31'b0010000000000010100001000000000,
31'b0010000000000100100001000000000,
31'b1010000010000000010000010000000,
31'b0010000000001000100001000000000,
31'b0010000000001010100001000000000,
31'b0010000000001100100001000000000,
31'b1100000000000001000000011000000,
31'b0001000000010000000110000000000,
31'b0010100000000000000011001000000,
31'b1001000000000000000000000110100,
31'b1000001010000000001000000000100,
31'b0001000010000000000000010010010,
31'b1100010010000000000000010000000,
31'b0100010000000000110001000000000,
31'b0100001001000001000000000000000,
31'b0001000000000000000110000000000,
31'b0001000000000010000110000000000,
31'b0100000000000001100000000100000,
31'b0100010000001000000100000000001,
31'b0001000000001000000110000000000,
31'b0101000010000001000000100000000,
31'b0100010000000010000100000000001,
31'b0100010000000000000100000000001,
31'b1000000000000000001100000010000,
31'b0000010000100000000000000100000,
31'b1000010000000000000001100000100,
31'b0000010000100100000000000100000,
31'b1000010000000000100000011000000,
31'b0010000000000001000000001010000,
31'b1000100000000000001000010000100,
31'b0110000000010000010000000100000,
31'b1000010101000000000010000000000,
31'b0000010000110000000000000100000,
31'b0000000100000010000001000010000,
31'b0000000100000000000001000010000,
31'b0100010100000010000000001000000,
31'b0100010100000000000000001000000,
31'b0110000000000010010000000100000,
31'b0110000000000000010000000100000,
31'b0000010000000010000000000100000,
31'b0000010000000000000000000100000,
31'b0000010000000110000000000100000,
31'b0000010000000100000000000100000,
31'b0000010000001010000000000100000,
31'b0000010000001000000000000100000,
31'b0101000000000000000010000100001,
31'b0100000110000001000000000000000,
31'b0000010000010010000000000100000,
31'b0000010000010000000000000100000,
31'b0000010001000000001000100010000,
31'b0000010000010100000000000100000,
31'b0000011001000000100000000000000,
31'b0000000000000001010001000000000,
31'b1010101000000000010000000000000,
31'b0010010010000000000000000010000,
31'b1000010100010000000010000000000,
31'b0000010001100000000000000100000,
31'b0110001000000000110000000000000,
31'b1000000100100000001000000000100,
31'b0001000100010000000001000001000,
31'b0010100000000000000000100100010,
31'b0001000000000000100000010000001,
31'b1001000000000000001100000001000,
31'b1000010100000000000010000000000,
31'b1000010100000010000010000000000,
31'b1000010100000100000010000000000,
31'b1000000000000000000100100100000,
31'b0001000100000000000001000001000,
31'b0101000000000000111000000000000,
31'b0001000100000100000001000001000,
31'b1101000100000000000000000000001,
31'b0000010001000010000000000100000,
31'b0000010001000000000000000100000,
31'b1000000100000010001000000000100,
31'b1000000100000000001000000000100,
31'b0000011000010000100000000000000,
31'b0000010001001000000000000100000,
31'b0001010000000000000000000111000,
31'b1100000000000000000000000101010,
31'b0000000000000000000101000000100,
31'b0000010001010000000000000100000,
31'b0000010000000000001000100010000,
31'b1000000100010000001000000000100,
31'b0000011000000000100000000000000,
31'b0000011000000010100000000000000,
31'b0000100000000000000001010010000,
31'b0010010011000000000000000010000,
31'b0100000000000010010000000010000,
31'b0100000000000000010000000010000,
31'b0100100001000001000000010000000,
31'b0100000000000100010000000010000,
31'b0100100100000000000000000001100,
31'b0100000000001000010000000010000,
31'b0101000001000000010000000001000,
31'b0100000100100001000000000000000,
31'b0100100000000000000000101000001,
31'b0100000000010000010000000010000,
31'b0000000000000011000000001100000,
31'b0000000000000001000000001100000,
31'b1001000001000000100100000000000,
31'b0100010110000000000000001000000,
31'b1010000000000000001100000100000,
31'b0010010000100000000000000010000,
31'b0101100000000000000100000000000,
31'b0000010010000000000000000100000,
31'b0101100000000100000100000000000,
31'b0100000100001001000000000000000,
31'b0101100000001000000100000000000,
31'b0100000100000101000000000000000,
31'b0100000100000011000000000000000,
31'b0100000100000001000000000000000,
31'b0110000000000010000001001000000,
31'b0110000000000000000001001000000,
31'b1010000000000000000000001001001,
31'b0010010000001000000000000010000,
31'b1010000001000000000011000000000,
31'b0010010000000100000000000010000,
31'b1000000000000001100000010000000,
31'b0010010000000000000000000010000,
31'b0100100000000101000000010000000,
31'b0100000001000000010000000010000,
31'b0100100000000001000000010000000,
31'b0100100000000011000000010000000,
31'b1001000000010000100100000000000,
31'b1010000000000000000100100010000,
31'b0101000000000000010000000001000,
31'b0101000000000010010000000001000,
31'b1001000000001000100100000000000,
31'b0100000001010000010000000010000,
31'b0100100000010001000000010000000,
31'b0000100000000000000000100010010,
31'b1001000000000000100100000000000,
31'b1001000000000010100100000000000,
31'b1100000000000001000010000100000,
31'b0010010001100000000000000010000,
31'b0101100001000000000100000000000,
31'b0100000000000000000000010001100,
31'b1000000100000001000010001000000,
31'b1000001000000001000000010100000,
31'b1010000000010000000011000000000,
31'b0100000101000101000000000000000,
31'b0101000000100000010000000001000,
31'b0100000101000001000000000000000,
31'b0011010000000000000000000001000,
31'b0110000001000000000001001000000,
31'b0011010000000100000000000001000,
31'b0011000000000000000010001000010,
31'b1010000000000000000011000000000,
31'b1010000000000010000011000000000,
31'b1010000000000100000011000000000,
31'b0010010001000000000000000010000,
31'b1000010001010000000010000000000,
31'b0000010100100000000000000100000,
31'b0000000000100000000110100000000,
31'b0000000000010000000001000010000,
31'b0100100010000000000000000001100,
31'b0100010000010000000000001000000,
31'b0100000010100011000000000000000,
31'b0100000010100001000000000000000,
31'b1000010001000000000010000000000,
31'b0000000000000100000001000010000,
31'b0000000000000010000001000010000,
31'b0000000000000000000001000010000,
31'b0100010000000010000000001000000,
31'b0100010000000000000000001000000,
31'b0100000000000000000010000001010,
31'b0000000000001000000001000010000,
31'b0000010100000010000000000100000,
31'b0000010100000000000000000100000,
31'b0000000000000000000110100000000,
31'b0010000000000000010000001000000,
31'b0100110000000000100010000000000,
31'b0100000010000101000000000000000,
31'b0100000010000011000000000000000,
31'b0100000010000001000000000000000,
31'b1000010001100000000010000000000,
31'b0000010100010000000000000100000,
31'b0000000000100010000001000010000,
31'b0000000000100000000001000010000,
31'b0100010000100010000000001000000,
31'b0100010000100000000000001000000,
31'b0100000010010011000000000000000,
31'b0100000010010001000000000000000,
31'b1000010000010000000010000000000,
31'b1000010000010010000010000000000,
31'b1000010000010100000010000000000,
31'b1000000000100000001000000000100,
31'b0001000000010000000001000001000,
31'b0101000010000000000100010000000,
31'b0001000100000000100000010000001,
31'b1101000000010000000000000000001,
31'b1000010000000000000010000000000,
31'b1000010000000010000010000000000,
31'b1000010000000100000010000000000,
31'b0000000001000000000001000010000,
31'b0001000000000000000001000001000,
31'b0100010001000000000000001000000,
31'b0001000000000100000001000001000,
31'b1101000000000000000000000000001,
31'b1000010000110000000010000000000,
31'b1000000000000100001000000000100,
31'b1000000000000010001000000000100,
31'b1000000000000000001000000000100,
31'b0001001000000000000000010010010,
31'b1100011000000000000000010000000,
31'b1110000000000000010010000000000,
31'b1000000000001000001000000000100,
31'b1000010000100000000010000000000,
31'b1000010000100010000010000000000,
31'b1000010000100100000010000000000,
31'b1000000000010000001000000000100,
31'b0001000000100000000001000001000,
31'b0101001000000001000000100000000,
31'b0001101000000000000000000100001,
31'b1101000000100000000000000000001,
31'b0100100000001000000000000001100,
31'b0100000100000000010000000010000,
31'b0100000000101011000000000000000,
31'b0100000000101001000000000000000,
31'b0100100000000000000000000001100,
31'b0010000000000000000001000100000,
31'b0100000000100011000000000000000,
31'b0100000000100001000000000000000,
31'b1000010011000000000010000000000,
31'b0010010000000001010000000000000,
31'b0000001000000001000010010000000,
31'b0000000010000000000001000010000,
31'b0100100000010000000000000001100,
31'b0100010010000000000000001000000,
31'b0100000010000000000010000001010,
31'b0100000000110001000000000000000,
31'b0101100100000000000100000000000,
31'b0100000000001101000000000000000,
31'b0100000000001011000000000000000,
31'b0100000000001001000000000000000,
31'b0100000000000111000000000000000,
31'b0100000000000101000000000000000,
31'b0100000000000011000000000000000,
31'b0100000000000001000000000000000,
31'b1000000001000000100000000001100,
31'b0110000100000000000001001000000,
31'b0100001000000000000101000000010,
31'b0100000000011001000000000000000,
31'b0100100000000000001000001000010,
31'b0100000000010101000000000000000,
31'b0100000000010011000000000000000,
31'b0100000000010001000000000000000,
31'b1000010010010000000010000000000,
31'b0101000000001000000100010000000,
31'b1000110000000000000000000000110,
31'b1000100000010001100000000000000,
31'b0101000000000010000100010000000,
31'b0101000000000000000100010000000,
31'b0101000100000000010000000001000,
31'b0100000001100001000000000000000,
31'b1000010010000000000010000000000,
31'b1000100000000101100000000000000,
31'b1000100000000011100000000000000,
31'b1000100000000001100000000000000,
31'b0010010000000000000100000000100,
31'b0101000000010000000100010000000,
31'b0010010000000100000100000000100,
31'b1101000010000000000000000000001,
31'b1000000000010000100000000001100,
31'b1000010000000001000000000001010,
31'b1000000000000001000010001000000,
31'b1000000010000000001000000000100,
31'b0100100000000000010000010010000,
31'b0100000001000101000000000000000,
31'b0100000001000011000000000000000,
31'b0100000001000001000000000000000,
31'b1000000000000000100000000001100,
31'b1000100000000000001010000000010,
31'b1000000000010001000010001000000,
31'b1000100000100001100000000000000,
31'b1010000100000000000011000000000,
31'b0100000001010101000000000000000,
31'b0100000001010011000000000000000,
31'b0100000001010001000000000000000,
31'b1101000000000000000000000000000,
31'b0000010000000000000000000010010,
31'b1101000000000100000000000000000,
31'b0001000000000000000001000001001,
31'b1101000000001000000000000000000,
31'b0001000001000000000010001000000,
31'b1101000000001100000000000000000,
31'b1000010000000000000010000000001,
31'b1101000000010000000000000000000,
31'b0001000100000000100000010000000,
31'b1101000000010100000000000000000,
31'b0001000100000100100000010000000,
31'b1101000000011000000000000000000,
31'b0001000100001000100000010000000,
31'b0010100000100000001000000100000,
31'b1110001000000000001000000000000,
31'b1101000000100000000000000000000,
31'b0001101000000000000000000100000,
31'b1101000000100100000000000000000,
31'b0001101000000100000000000100000,
31'b1101000000101000000000000000000,
31'b0010100001000000000000100010000,
31'b0010100000010000001000000100000,
31'b1100000000000000010000010000100,
31'b1101000000110000000000000000000,
31'b0001101000010000000000000100000,
31'b0010100000001000001000000100000,
31'b0000100000000000100000000011000,
31'b1000000000000000001000000000101,
31'b1001001000000000000010010000000,
31'b0010100000000000001000000100000,
31'b0110000000000000010000000010010,
31'b1101000001000000000000000000000,
31'b0001000000001000000010001000000,
31'b1000000000000000000011000000010,
31'b1100000000001000000000000011000,
31'b0000000000000000000001000010001,
31'b0001000000000000000010001000000,
31'b0001010000000000000000000001010,
31'b1100000000000000000000000011000,
31'b1101000001010000000000000000000,
31'b0001000101000000100000010000000,
31'b1100001010000000000000100000000,
31'b0010001010000001000000000000100,
31'b0001100000100000100000000000000,
31'b0001000000010000000010001000000,
31'b0001100000100100100000000000000,
31'b1100000000010000000000000011000,
31'b1101000001100000000000000000000,
31'b0010100000001000000000100010000,
31'b1100000000000001000100010000000,
31'b0010101000000000101000000000000,
31'b0001100000010000100000000000000,
31'b0010100000000000000000100010000,
31'b0001100000010100100000000000000,
31'b1100000000100000000000000011000,
31'b0100000010000001000000000000001,
31'b0101000100000000000010000100000,
31'b0101010000000000000100100000000,
31'b0000100010000000000000100100000,
31'b0001100000000000100000000000000,
31'b0001100000000010100000000000000,
31'b0001100000000100100000000000000,
31'b0001100000000110100000000000000,
31'b1101000010000000000000000000000,
31'b0001000000000000011100000000000,
31'b1101000010000100000000000000000,
31'b0010010000000000000100000000101,
31'b1101000010001000000000000000000,
31'b0001000011000000000010001000000,
31'b0010001000010000010100000000000,
31'b1100000000000000100000100100000,
31'b1101000010010000000000000000000,
31'b0001000110000000100000010000000,
31'b1100001001000000000000100000000,
31'b0010010000001000000000000100010,
31'b0010001000000100010100000000000,
31'b0000010000000000000110010000000,
31'b0010001000000000010100000000000,
31'b0010010000000000000000000100010,
31'b0000100000000000001000000010000,
31'b0100000000000000010000000100010,
31'b0100000000000000000000111000000,
31'b0100000000000100010000000100010,
31'b0100000000000000100001000000100,
31'b0100000000001000010000000100010,
31'b0000101000000000100000100000000,
31'b1000000001000000000010110000000,
31'b0100000001000001000000000000001,
31'b0100000001000011000000000000001,
31'b0100000001000101000000000000001,
31'b0000100001000000000000100100000,
31'b1001000000000001000001000010000,
31'b1000000100000000000001010000100,
31'b0010100010000000001000000100000,
31'b0011101000000000000000000010000,
31'b1101000011000000000000000000000,
31'b0001000010001000000010001000000,
31'b1100001000010000000000100000000,
31'b0010001000010001000000000000100,
31'b0001000000000001001000000000100,
31'b0001000010000000000010001000000,
31'b0010010000000001010000000000001,
31'b1100000010000000000000000011000,
31'b1000100000000000000001000000100,
31'b1110000000000000000000000101000,
31'b1100001000000000000000100000000,
31'b0010001000000001000000000000100,
31'b1100000000000000101000000010000,
31'b0001010000000000101000000000010,
31'b1100001000001000000000100000000,
31'b0010010001000000000000000100010,
31'b0100000000010001000000000000001,
31'b0100000001000000010000000100010,
31'b0100000001000000000000111000000,
31'b0000100000010000000000100100000,
31'b0100000001000000100001000000100,
31'b1010000100000000000000001001000,
31'b1000001000000000000100000001010,
31'b1000000000000000000010110000000,
31'b0100000000000001000000000000001,
31'b0100000000000011000000000000001,
31'b0100000000000101000000000000001,
31'b0000100000000000000000100100000,
31'b0100000000001001000000000000001,
31'b0100010000000000100100000100000,
31'b0100000100000000100010100000000,
31'b0001010000000001000010000000000,
31'b1101000100000000000000000000000,
31'b0001000000010000100000010000000,
31'b1101000100000100000000000000000,
31'b0001000100000000000001000001001,
31'b1101000100001000000000000000000,
31'b0001000101000000000010001000000,
31'b0010100000000000000100100000100,
31'b1100100000000001000100000000000,
31'b1000000000000000000000100000110,
31'b0001000000000000100000010000000,
31'b1001000010000000010001000000000,
31'b0001000000000100100000010000000,
31'b1001000000100000000000001100000,
31'b0001000000001000100000010000000,
31'b0000000010000000000000110100000,
31'b0001000000001100100000010000000,
31'b1101000100100000000000000000000,
31'b0001101100000000000000000100000,
31'b0000011000000010100000000000001,
31'b0000011000000000100000000000001,
31'b1100000000000000000100000001100,
31'b0010000010000000000001000010010,
31'b0000001000000001000100000100000,
31'b0000010000000001010000000000010,
31'b1001000000001000000000001100000,
31'b0001000000100000100000010000000,
31'b0000000000001000110000000000100,
31'b0000000000000000000001000100010,
31'b1001000000000000000000001100000,
31'b1001000000000010000000001100000,
31'b0000000000000000110000000000100,
31'b0000000000001000000001000100010,
31'b1101000101000000000000000000000,
31'b0001000100001000000010001000000,
31'b1100100000000000010000000000100,
31'b0010100000000001010000100000000,
31'b0001001000000000000000010100000,
31'b0001000100000000000010001000000,
31'b0001010100000000000000000001010,
31'b1100000100000000000000000011000,
31'b1001101000000000000010000000000,
31'b0001000001000000100000010000000,
31'b0010000000000010001000010100000,
31'b0010000000000000001000010100000,
31'b0001100100100000100000000000000,
31'b0001000100010000000010001000000,
31'b0000010000100000000000000100001,
31'b1010010000000001000000000001000,
31'b0010010010000000000000000010001,
31'b1100000000000001010000000001000,
31'b0000010000000000000100000000110,
31'b0000001000000000010000000100100,
31'b0001100100010000100000000000000,
31'b1101100000000000000000010000000,
31'b0000010000010000000000000100001,
31'b0000010001000001010000000000010,
31'b0101000000000010000010000100000,
31'b0101000000000000000010000100000,
31'b0000010000001000000000000100001,
31'b0000000000000001100100000000000,
31'b0001100100000000100000000000000,
31'b0101000000001000000010000100000,
31'b0000010000000000000000000100001,
31'b0000010000000010000000000100001,
31'b1101000110000000000000000000000,
31'b0001000100000000011100000000000,
31'b1000100000000000000010100000000,
31'b1001000000000000100100000000001,
31'b0000100000000101011000000000000,
31'b0000000001000000001000010010000,
31'b0000100000000001011000000000000,
31'b0100100001000000000000101000000,
31'b1001000000000100010001000000000,
31'b0001000010000000100000010000000,
31'b1001000000000000010001000000000,
31'b1001000000000010010001000000000,
31'b0000000000000100000000110100000,
31'b0000000000000000010000001000010,
31'b0000000000000000000000110100000,
31'b0000000000000100010000001000010,
31'b0110000000000000000010000001000,
31'b0110000000000010000010000001000,
31'b1011000000000000000000001010000,
31'b1010000000000000000011000000001,
31'b0110000000001000000010000001000,
31'b0010000000000000000001000010010,
31'b0000101100000000100000100000000,
31'b0011010000000000000000000001001,
31'b0110000000010000000010000001000,
31'b1000000000001000000001010000100,
31'b1001000000100000010001000000000,
31'b1000000000000000100000101000000,
31'b1001000010000000000000001100000,
31'b1000000000000000000001010000100,
31'b0000000010000000110000000000100,
31'b1000000000001000100000101000000,
31'b0010010000100000000000000010001,
31'b0000010000000000100100001000000,
31'b1001001000000000000000000000110,
31'b0000100000000000001100000000100,
31'b0000000000000010001000010010000,
31'b0000000000000000001000010010000,
31'b0100100000000010000000101000000,
31'b0100100000000000000000101000000,
31'b1100000000000000010010000000010,
31'b0001010000000000010010000010000,
31'b1100001100000000000000100000000,
31'b0010001100000001000000000000100,
31'b0100000000000100010000000010001,
31'b0000000001000000010000001000010,
31'b0100000000000000010000000010001,
31'b0100100000010000000000101000000,
31'b0010010000000000000000000010001,
31'b1010000000001000000000001001000,
31'b0011000000000000000001000001010,
31'b0000100100010000000000100100000,
31'b1010000000000010000000001001000,
31'b1010000000000000000000001001000,
31'b1010010000000000000010000000010,
31'b1010000000000100000000001001000,
31'b0100000100000001000000000000001,
31'b0101000010000000000010000100000,
31'b0100000100000101000000000000001,
31'b0000100100000000000000100100000,
31'b0100000100001001000000000000001,
31'b1010000000010000000000001001000,
31'b0100000000000000100010100000000,
31'b0101100000000000000100000000001,
31'b1101001000000000000000000000000,
31'b0001100000100000000000000100000,
31'b1101001000000100000000000000000,
31'b0001100000100100000000000100000,
31'b1101001000001000000000000000000,
31'b0001100000101000000000000100000,
31'b0010000100000000101000010000000,
31'b1110000000010000001000000000000,
31'b1101001000010000000000000000000,
31'b0001100000110000000000000100000,
31'b1000000000000000010010000000100,
31'b1110000000001000001000000000000,
31'b0010000010000100010100000000000,
31'b1110000000000100001000000000000,
31'b0010000010000000010100000000000,
31'b1110000000000000001000000000000,
31'b0100010010000000000100000000000,
31'b0001100000000000000000000100000,
31'b0101000000000001000000100000001,
31'b0001100000000100000000000100000,
31'b0101000100000000100010000000000,
31'b0001100000001000000000000100000,
31'b0000100010000000100000100000000,
31'b0001100000001100000000000100000,
31'b0101000001000000000000011000000,
31'b0001100000010000000000000100000,
31'b1100010000000000000000010000001,
31'b0001100000010100000000000100000,
31'b1001000000000010000010010000000,
31'b1001000000000000000010010000000,
31'b0010101000000000001000000100000,
31'b1110000000100000001000000000000,
31'b1101001001000000000000000000000,
31'b0010100000000001000010000000010,
31'b1100000010010000000000100000000,
31'b0010100000100000101000000000000,
31'b0001000100000000000000010100000,
31'b0001001000000000000010001000000,
31'b0001011000000000000000000001010,
31'b1100001000000000000000000011000,
31'b1100000010000100000000100000000,
31'b0010010000000000001000000001010,
31'b1100000010000000000000100000000,
31'b0010000010000001000000000000100,
31'b0001101000100000100000000000000,
31'b1101000000000000100000000100000,
31'b1100000010001000000000100000000,
31'b1000000000000001000110000000000,
31'b0101000000010000000000011000000,
31'b0010010000000000000000001000100,
31'b0010100000000010101000000000000,
31'b0010100000000000101000000000000,
31'b0001101000010000100000000000000,
31'b0010101000000000000000100010000,
31'b0000100000000000000000000111000,
31'b0110000000000000000001000010100,
31'b0101000000000000000000011000000,
31'b0101000000000010000000011000000,
31'b1100000010100000000000100000000,
31'b0010100000010000101000000000000,
31'b0001101000000000100000000000000,
31'b1001000001000000000010010000000,
31'b0001101000000100100000000000000,
31'b1100000000000000000001010000010,
31'b1000100000000000010000000000010,
31'b1100000000000000001000000110000,
31'b1100000001010000000000100000000,
31'b0010000001010001000000000000100,
31'b1110000000000000100000000001000,
31'b0010000100010000000000010001000,
31'b0010000000010000010100000000000,
31'b0010000000000000100001000000001,
31'b1100000001000100000000100000000,
31'b0010000100001000000000010001000,
31'b1100000001000000000000100000000,
31'b0010000001000001000000000000100,
31'b0010000000000100010100000000000,
31'b0010000100000000000000010001000,
31'b0010000000000000010100000000000,
31'b0000000000000000000010101000000,
31'b0100010000000000000100000000000,
31'b0100010000000010000100000000000,
31'b0100010000000100000100000000000,
31'b0100010000000110000100000000000,
31'b0100010000001000000100000000000,
31'b0100010000001010000100000000000,
31'b0000100000000000100000100000000,
31'b0001000000000000000110000000001,
31'b0100010000010000000100000000000,
31'b0100010000010010000100000000000,
31'b1100000001100000000000100000000,
31'b0011100000001000000000000010000,
31'b0100010000011000000100000000000,
31'b1001000010000000000010010000000,
31'b0010000000100000010100000000000,
31'b0011100000000000000000000010000,
31'b1100000000010100000000100000000,
31'b0010000000010101000000000000100,
31'b1100000000010000000000100000000,
31'b0010000000010001000000000000100,
31'b0001001000000001001000000000100,
31'b0000000100000000000001001000100,
31'b1100000000011000000000100000000,
31'b0010000001000000100001000000001,
31'b1100000000000100000000100000000,
31'b0010000000000101000000000000100,
31'b1100000000000000000000100000000,
31'b0010000000000001000000000000100,
31'b1100000000001100000000100000000,
31'b0010000101000000000000010001000,
31'b1100000000001000000000100000000,
31'b0010000000001001000000000000100,
31'b0100010001000000000100000000000,
31'b0100010001000010000100000000000,
31'b1100000000110000000000100000000,
31'b0010100010000000101000000000000,
31'b1010010000000000010000100000000,
31'b1000010000000000000110001000000,
31'b1000000000000000000100000001010,
31'b1000001000000000000010110000000,
31'b0010100000000000000000000001000,
31'b0100000000000000000001000100100,
31'b1100000000100000000000100000000,
31'b0010000000100001000000000000100,
31'b0100000000000000110000000000010,
31'b0100000000001000000001000100100,
31'b1100000000101000000000100000000,
31'b0011100001000000000000000010000,
31'b1101001100000000000000000000000,
31'b0001100100100000000000000100000,
31'b0010010000000000000100001010000,
31'b0000010000100000100000000000001,
31'b0110000000000000000101000000000,
31'b0110000000000010000101000000000,
31'b0010000000000000101000010000000,
31'b1010000000000000000100000001001,
31'b1001100001000000000010000000000,
31'b0001001000000000100000010000000,
31'b1100100000000000000001000000010,
31'b0001110000000000000001000010000,
31'b0110000000010000000101000000000,
31'b0101100000000000000000001000000,
31'b0010000110000000010100000000000,
31'b1110000100000000001000000000000,
31'b0101000000001000100010000000000,
31'b0001100100000000000000000100000,
31'b0000010000000010100000000000001,
31'b0000010000000000100000000000001,
31'b0101000000000000100010000000000,
31'b0101000000000010100010000000000,
31'b0000000000000001000100000100000,
31'b0000010000001000100000000000001,
31'b0010000010000001000100000010000,
31'b0001100100010000000000000100000,
31'b0000010000000000010101000000000,
31'b0000010000010000100000000000001,
31'b1001001000000000000000001100000,
31'b1001000100000000000010010000000,
31'b0000001000000000110000000000100,
31'b0000010001000001000001000000100,
31'b1000000000000000010001100000000,
31'b1001000000100000100000001000000,
31'b1001000010000000000000000000110,
31'b0000000010000000100000110000000,
31'b0001000000000000000000010100000,
31'b0001000000000010000000010100000,
31'b0001000000000100000000010100000,
31'b0001000000000110000000010100000,
31'b1001100000000000000010000000000,
31'b1001100000000010000010000000000,
31'b1100000110000000000000100000000,
31'b0010001000000000001000010100000,
31'b0001000000010000000000010100000,
31'b0110010000000000000000000100100,
31'b0001100000000000000000000010011,
31'b1100110000000000000000000000001,
31'b1001000000000010100000001000000,
31'b1001000000000000100000001000000,
31'b0000000000001000100001000000010,
31'b0000000000000000010000000100100,
31'b0001000000100000000000010100000,
31'b1001000000001000100000001000000,
31'b0000000000000000100001000000010,
31'b0000000000001000010000000100100,
31'b1010000000000000000000101010000,
31'b1001000000010000100000001000000,
31'b0000011000001000000000000100001,
31'b0000001000000001100100000000000,
31'b0001101100000000100000000000000,
31'b0010010000000000000000100001001,
31'b0000011000000000000000000100001,
31'b0000010000000001000001000000100,
31'b1100000000000000000011000000100,
31'b0010000000011000000000010001000,
31'b1001000001000000000000000000110,
31'b0000000001000000100000110000000,
31'b0110000010000000000101000000000,
31'b0010000000010000000000010001000,
31'b0010000100010000010100000000000,
31'b0010000100000000100001000000001,
31'b0010000000100001000100000010000,
31'b0010000000001000000000010001000,
31'b1100000101000000000000100000000,
31'b0010000101000001000000000000100,
31'b0010000000000010000000010001000,
31'b0010000000000000000000010001000,
31'b0010000100000000010100000000000,
31'b0010000000000100000000010001000,
31'b0100010100000000000100000000000,
31'b0100010100000010000100000000000,
31'b0100010100000100000100000000000,
31'b0100000000000000000010100100000,
31'b0101000010000000100010000000000,
31'b1000000001000000010000010000010,
31'b0000100100000000100000100000000,
31'b0101110000000001000000000000000,
31'b0010000000000001000100000010000,
31'b1000010000000000100100010000000,
31'b0011000000000000010000000001100,
31'b1100010000000000001001000000000,
31'b1000000000000010001000001010000,
31'b1000000000000000001000001010000,
31'b0010100000000001000000010000100,
31'b1100100000000000000000110000000,
31'b1001000000000100000000000000110,
31'b0000000000001000000001001000100,
31'b1001000000000000000000000000110,
31'b0000000000000000100000110000000,
31'b0001000010000000000000010100000,
31'b0000000000000000000001001000100,
31'b1001000000001000000000000000110,
31'b0000000000001000100000110000000,
31'b1100000100000100000000100000000,
31'b0010000100000101000000000000100,
31'b1100000100000000000000100000000,
31'b0010000100000001000000000000100,
31'b0011100000000000000100000000100,
31'b0010000001000000000000010001000,
31'b1100000100001000000000100000000,
31'b0010000100001001000000000000100,
31'b0100010101000000000100000000000,
31'b1001000010000000100000001000000,
31'b1001000000100000000000000000110,
31'b0000000010000000010000000100100,
31'b1000000000000100000000101100000,
31'b1000000000000000010000010000010,
31'b1000000000000000000000101100000,
31'b1000000000000100010000010000010,
31'b0100000000000000001010000010000,
31'b0100000100000000000001000100100,
31'b1100000100100000000000100000000,
31'b0010100000000000010100010000000,
31'b0100000100000000110000000000010,
31'b0010000000000000010000000010100,
31'b1100000000000000001000000000011,
31'b0011000000000001000100000001000,
31'b0000000000000010000000000010010,
31'b0000000000000000000000000010010,
31'b0100000001000000000000001000001,
31'b0000000000000100000000000010010,
31'b0100000000000000000011000001000,
31'b0000000000001000000000000010010,
31'b1000000000000010000010000000001,
31'b1000000000000000000010000000001,
31'b0100000000000001000000110000000,
31'b0000000000010000000000000010010,
31'b0100000001010000000000001000001,
31'b0000100000000000000000010100001,
31'b0100000000010000000011000001000,
31'b0000000010000000000110010000000,
31'b1011000000100000010000000000000,
31'b1000000000010000000010000000001,
31'b0100001010000000000100000000000,
31'b0000000000100000000000000010010,
31'b0100001010000100000100000000000,
31'b0000001100000000100000000000001,
31'b0100001010001000000100000000000,
31'b0000001000000001000010100000000,
31'b1011000000010000010000000000000,
31'b1000000000100000000010000000001,
31'b0100001010010000000100000000000,
31'b0000001000000000000001010001000,
31'b1100001000000000000000010000001,
31'b0000110000000000100000000011000,
31'b1011000000000100010000000000000,
31'b0100000010000001000001000000010,
31'b1011000000000000010000000000000,
31'b1011000000000010010000000000000,
31'b0100000000000100000000001000001,
31'b0000000001000000000000000010010,
31'b0100000000000000000000001000001,
31'b0100000000000010000000001000001,
31'b0001000000000100000000000001010,
31'b0001010000000000000010001000000,
31'b0001000000000000000000000001010,
31'b1000000001000000000010000000001,
31'b0100000001000001000000110000000,
31'b0000000001010000000000000010010,
31'b0100000000010000000000001000001,
31'b0100100000000000010000100010000,
31'b0001110000100000100000000000000,
31'b0001010000010000000010001000000,
31'b0001000000010000000000000001010,
31'b1010000100000001000000000001000,
31'b0100001011000000000100000000000,
31'b0010001000000000000000001000100,
31'b0100000000100000000000001000001,
31'b0110000000000000100100000010000,
31'b0001110000010000100000000000000,
31'b0010110000000000000000100010000,
31'b0001000000100000000000000001010,
31'b1000000010000000010000000101000,
31'b0101000000000100000100100000000,
31'b1010000000000000010000000011000,
31'b0101000000000000000100100000000,
31'b0101000000000010000100100000000,
31'b0001110000000000100000000000000,
31'b0100100100000001000000100000000,
31'b0000000100000000000000000100001,
31'b0001000010000001000010000000000,
31'b0100001000100000000100000000000,
31'b0000000010000000000000000010010,
31'b0100001000100100000100000000000,
31'b0010000000000000000100000000101,
31'b0100001000101000000100000000000,
31'b0000000010001000000000000010010,
31'b1001000100000001000000000100000,
31'b1000000010000000000010000000001,
31'b0100001000110000000100000000000,
31'b0000000010010000000000000010010,
31'b0010000000001010000000000100010,
31'b0010000000001000000000000100010,
31'b0000001000000000000000100001010,
31'b0000000000000000000110010000000,
31'b0010000000000010000000000100010,
31'b0010000000000000000000000100010,
31'b0100001000000000000100000000000,
31'b0100001000000010000100000000000,
31'b0100001000000100000100000000000,
31'b0110000100000000000000001000010,
31'b0100001000001000000100000000000,
31'b0100001000001010000100000000000,
31'b0100100000000000001001001000000,
31'b1000000010100000000010000000001,
31'b0100001000010000000100000000000,
31'b0100001000010010000100000000000,
31'b1101000000000001000000001000000,
31'b0011000000000000000000101000100,
31'b0100001000011000000100000000000,
31'b0100000000000001000001000000010,
31'b1011000010000000010000000000000,
31'b0010000000100000000000000100010,
31'b0100001001100000000100000000000,
31'b0000000100000000100100001000000,
31'b0100000010000000000000001000001,
31'b0100001100000000000000000010100,
31'b0010000000000101010000000000001,
31'b0001010010000000000010001000000,
31'b0010000000000001010000000000001,
31'b1000000011000000000010000000001,
31'b1100000000000000000100011000000,
31'b0001000100000000010010000010000,
31'b1100011000000000000000100000000,
31'b0010011000000001000000000000100,
31'b1000101000000000100100000000000,
31'b0001000000000000101000000000010,
31'b0010000001000010000000000100010,
31'b0010000001000000000000000100010,
31'b0100001001000000000100000000000,
31'b0100001001000010000100000000000,
31'b0100001001000100000100000000000,
31'b1000100000000000001011000000000,
31'b1010001000000000010000100000000,
31'b1000001000000000000110001000000,
31'b1010000100000000000010000000010,
31'b1000000000000000010000000101000,
31'b0100010000000001000000000000001,
31'b0100010000000011000000000000001,
31'b0101000010000000000100100000000,
31'b0001000000001001000010000000000,
31'b0100010000001001000000000000001,
31'b0100000000000000100100000100000,
31'b0001000000000011000010000000000,
31'b0001000000000001000010000000000,
31'b0110000000000000100000000000100,
31'b0000000100000000000000000010010,
31'b0110000000000100100000000000100,
31'b0000001000100000100000000000001,
31'b0110000000001000100000000000100,
31'b0000000100001000000000000010010,
31'b1001000010000001000000000100000,
31'b1000000100000000000010000000001,
31'b1011000000000001000000000010000,
31'b0001010000000000100000010000000,
31'b0000101000000000000010001000001,
31'b0001101000000000000001000010000,
31'b0000101001000000000001000001000,
31'b0001010000001000100000010000000,
31'b0000000010000000010010000001000,
31'b1010000001000001000000000001000,
31'b0110000000100000100000000000100,
31'b0000001000000100100000000000001,
31'b0000001000000010100000000000001,
31'b0000001000000000100000000000001,
31'b0000100001000000000000010010010,
31'b0000000000000101010000000000010,
31'b0000000001010000000000000100001,
31'b0000000000000001010000000000010,
31'b0000100011000000000110000000000,
31'b0001010000100000100000010000000,
31'b0000001000000000010101000000000,
31'b0000010000000000000001000100010,
31'b0000100000000000011000001000000,
31'b0100100001000001000000100000000,
31'b0000000001000000000000000100001,
31'b0000000001000010000000000100001,
31'b0110000001000000100000000000100,
31'b0000000101000000000000000010010,
31'b0100000100000000000000001000001,
31'b0100001010000000000000000010100,
31'b0001011000000000000000010100000,
31'b0001010100000000000010001000000,
31'b0001000100000000000000000001010,
31'b1010000000010001000000000001000,
31'b0000101000001000000001000001000,
31'b0001010001000000100000010000000,
31'b0000000000101000000000000100001,
31'b1010000000001001000000000001000,
31'b0000101000000000000001000001000,
31'b1010000000000101000000000001000,
31'b0000000000100000000000000100001,
31'b1010000000000001000000000001000,
31'b0010000010000000000000000010001,
31'b0010001100000000000000001000100,
31'b0000000000000000000100000000110,
31'b0000001001000000100000000000001,
31'b0000100000000000000000010010010,
31'b0100100000010001000000100000000,
31'b0000000000010000000000000100001,
31'b0000000001000001010000000000010,
31'b0000100010000000000110000000000,
31'b0101010000000000000010000100000,
31'b0000000000001000000000000100001,
31'b0000010000000001100100000000000,
31'b0000000000000100000000000100001,
31'b0100100000000001000000100000000,
31'b0000000000000000000000000100001,
31'b0000000000000010000000000100001,
31'b0110000010000000100000000000100,
31'b0000000110000000000000000010010,
31'b1001000000001001000000000100000,
31'b0110000000100000000000001000010,
31'b1100000000000000100110000000000,
31'b0000010001000000001000010010000,
31'b1001000000000001000000000100000,
31'b1001000000000011000000000100000,
31'b0000100001100000000110000000000,
31'b0001010010000000100000010000000,
31'b0000100000000000001001000100000,
31'b0110000000000000001000000001100,
31'b0000001000000000000100001100000,
31'b0000010000000000010000001000010,
31'b0000000000000000010010000001000,
31'b0010000100000000000000000100010,
31'b0100001100000000000100000000000,
31'b0110000000000100000000001000010,
31'b0110000000000010000000001000010,
31'b0110000000000000000000001000010,
31'b1111000000000000000001000000000,
31'b0011000000000100000000000001001,
31'b1010000001000000000010000000010,
31'b0011000000000000000000000001001,
31'b0000100001000000000110000000000,
31'b1000100000000000001000100000100,
31'b0000100001000100000110000000000,
31'b1100001000000000001001000000000,
31'b0000100010000000011000001000000,
31'b1100100000000000000100001000000,
31'b0000000011000000000000000100001,
31'b0011000000010000000000000001001,
31'b0010000000100000000000000010001,
31'b0000000000000000100100001000000,
31'b0100001000000010000000000010100,
31'b0100001000000000000000000010100,
31'b1010000000000001101000000000000,
31'b0000010000000000001000010010000,
31'b1010000000100000000010000000010,
31'b0100110000000000000000101000000,
31'b0000100000100000000110000000000,
31'b0001000000000000010010000010000,
31'b0000100001000000001001000100000,
31'b1100000000000000010000001001000,
31'b0000101010000000000001000001000,
31'b0001000100000000101000000000010,
31'b0000000010100000000000000100001,
31'b1010000010000001000000000001000,
31'b0010000000000000000000000010001,
31'b0010000000000010000000000010001,
31'b0010000000000100000000000010001,
31'b0110000001000000000000001000010,
31'b1000000000000000000100010100000,
31'b1010010000000000000000001001000,
31'b1010000000000000000010000000010,
31'b1010000000000010000010000000010,
31'b0000100000000000000110000000000,
31'b0001000000000000100000100000001,
31'b0000100000000100000110000000000,
31'b0001000100001001000010000000000,
31'b0000100000001000000110000000000,
31'b0100100010000001000000100000000,
31'b0000000010000000000000000100001,
31'b0001000100000001000010000000000,
31'b0100000010100000000100000000000,
31'b0000001000000000000000000010010,
31'b0100001001000000000000001000001,
31'b0000001000000100000000000010010,
31'b0100001000000000000011000001000,
31'b0000001000001000000000000010010,
31'b1001000000000000001000010000100,
31'b1000001000000000000010000000001,
31'b0100001000000001000000110000000,
31'b0000001000010000000000000010010,
31'b1100000000100000000000010000001,
31'b0001100100000000000001000010000,
31'b0000000010000000000000100001010,
31'b0000001010000000000110010000000,
31'b0011000000000000001000000010010,
31'b1110010000000000001000000000000,
31'b0100000010000000000100000000000,
31'b1000000000000000011000000000000,
31'b0100000010000100000100000000000,
31'b0000000100000000100000000000001,
31'b0100000010001000000100000000000,
31'b0000000000000001000010100000000,
31'b0100100000000000000010000100001,
31'b0000000100001000100000000000001,
31'b0100000010010000000100000000000,
31'b0000000000000000000001010001000,
31'b1100000000000000000000010000001,
31'b0000000100010000100000000000001,
31'b0100000010011000000100000000000,
31'b0000000000010001000010100000000,
31'b1100000000001000000000010000001,
31'b0000000101000001000001000000100,
31'b0100001000000100000000001000001,
31'b0010000000100000000000001000100,
31'b0100001000000000000000001000001,
31'b0100001000000010000000001000001,
31'b0001010100000000000000010100000,
31'b0011000000000000000000100100010,
31'b0001001000000000000000000001010,
31'b1000100000000000001100000001000,
31'b0010100000000000100010000000100,
31'b0010000000000000001000000001010,
31'b1100010010000000000000100000000,
31'b0010010010000001000000000000100,
31'b0000100100000000000001000001000,
31'b0110000100000000000000000100100,
31'b0001001000010000000000000001010,
31'b1100100100000000000000000000001,
31'b0100000011000000000100000000000,
31'b0010000000000000000000001000100,
31'b0100001000100000000000001000001,
31'b0010000000000100000000001000100,
31'b1010000010000000010000100000000,
31'b0010000000001000000000001000100,
31'b0001001000100000000000000001010,
31'b0010000000001100000000001000100,
31'b0101010000000000000000011000000,
31'b0010000000010000000000001000100,
31'b1100000001000000000000010000001,
31'b0010000000010100000000001000100,
31'b0001111000000000100000000000000,
31'b0010000100000000000000100001001,
31'b0001000000000000000001010010000,
31'b0000000100000001000001000000100,
31'b0100000000100000000100000000000,
31'b0100000000100010000100000000000,
31'b0100000000100100000100000000000,
31'b0100000101000000000000000010100,
31'b0100000000101000000100000000000,
31'b0100000000101010000100000000000,
31'b0100100001000000010000000001000,
31'b1000001010000000000010000000001,
31'b0100000000110000000100000000000,
31'b0100000000110010000100000000000,
31'b1100010001000000000000100000000,
31'b0010010001000001000000000000100,
31'b0000000000000000000000100001010,
31'b0000001000000000000110010000000,
31'b0010010000000000010100000000000,
31'b0010001000000000000000000100010,
31'b0100000000000000000100000000000,
31'b0100000000000010000100000000000,
31'b0100000000000100000100000000000,
31'b0100000000000110000100000000000,
31'b0100000000001000000100000000000,
31'b0100000000001010000100000000000,
31'b0100000000001100000100000000000,
31'b0101100100000001000000000000000,
31'b0100000000010000000100000000000,
31'b0100000000010010000100000000000,
31'b1000000000000000110000000001000,
31'b1100000100000000001001000000000,
31'b0100000000011000000100000000000,
31'b0100001000000001000001000000010,
31'b1110100000000000000000000000010,
31'b0011110000000000000000000010000,
31'b0100000001100000000100000000000,
31'b0100000100000100000000000010100,
31'b0010000000000000100000000000010,
31'b0100000100000000000000000010100,
31'b1010000000100000010000100000000,
31'b1000100000000000010001000000001,
31'b0100100000000000010000000001000,
31'b0100100000000010010000000001000,
31'b1100010000000100000000100000000,
31'b0010010000000101000000000000100,
31'b1100010000000000000000100000000,
31'b0010010000000001000000000000100,
31'b1000100000000000100100000000000,
31'b1001000000000000000010100000001,
31'b1100010000001000000000100000000,
31'b0010010000001001000000000000100,
31'b0100000001000000000100000000000,
31'b0100000001000010000100000000000,
31'b0100000001000100000100000000000,
31'b0100000100100000000000000010100,
31'b1010000000000000010000100000000,
31'b1000000000000000000110001000000,
31'b1010000000000100010000100000000,
31'b1000001000000000010000000101000,
31'b0100000001010000000100000000000,
31'b0100010000000000000001000100100,
31'b1100010000100000000000100000000,
31'b0010100000000000000010001000010,
31'b1010000000010000010000100000000,
31'b1001000000000000110000000010000,
31'b0001001000000011000010000000000,
31'b0001001000000001000010000000000,
31'b0110001000000000100000000000100,
31'b0000001100000000000000000010010,
31'b0010000000000000000100001010000,
31'b0000000000100000100000000000001,
31'b0110010000000000000101000000000,
31'b1000000000000101001000000010000,
31'b1000000000000011001000000010000,
31'b1000000000000001001000000010000,
31'b0000100001001000000001000001000,
31'b0001100000000100000001000010000,
31'b0000100000000000000010001000001,
31'b0001100000000000000001000010000,
31'b0000100001000000000001000001000,
31'b0110000001000000000000000100100,
31'b0000100001000100000001000001000,
31'b1100100001000000000000000000001,
31'b0100000110000000000100000000000,
31'b0000000000000100100000000000001,
31'b0000000000000010100000000000001,
31'b0000000000000000100000000000001,
31'b0101010000000000100010000000000,
31'b0000000100000001000010100000000,
31'b0000010000000001000100000100000,
31'b0000000000001000100000000000001,
31'b0000000010000000001000000001001,
31'b0000000100000000000001010001000,
31'b0000000000000000010101000000000,
31'b0000000000010000100000000000001,
31'b0000101000000000011000001000000,
31'b0010000001000000000000100001001,
31'b0000001001000000000000000100001,
31'b0000000001000001000001000000100,
31'b1001000000000001001000000001000,
31'b0110000000000000000100000000011,
31'b0100001100000000000000001000001,
31'b0100000010000000000000000010100,
31'b0001010000000000000000010100000,
31'b0110000000010000000000000100100,
31'b0001010000000100000000010100000,
31'b1100100000010000000000000000001,
31'b0000100000001000000001000001000,
31'b0110000000001000000000000100100,
31'b0000100001000000000010001000001,
31'b1100100000001000000000000000001,
31'b0000100000000000000001000001000,
31'b0110000000000000000000000100100,
31'b0000100000000100000001000001000,
31'b1100100000000000000000000000001,
31'b0100000111000000000100000000000,
31'b0010000100000000000000001000100,
31'b0000001000000000000100000000110,
31'b0000000001000000100000000000001,
31'b0001010000100000000000010100000,
31'b0010000100001000000000001000100,
31'b0000010000000000100001000000010,
31'b0000000001001000100000000000001,
31'b0000101010000000000110000000000,
31'b0010000100010000000000001000100,
31'b0000001000001000000000000100001,
31'b0000000001010000100000000000001,
31'b0000100000100000000001000001000,
31'b0010000000000000000000100001001,
31'b0000001000000000000000000100001,
31'b0000000000000001000001000000100,
31'b0100000100100000000100000000000,
31'b0100000100100010000100000000000,
31'b0100000100100100000100000000000,
31'b0100000001000000000000000010100,
31'b0101000000000000000000000001100,
31'b0101000000000010000000000001100,
31'b1001001000000001000000000100000,
31'b1001000000000000000001000000101,
31'b0000000000100000001000000001001,
31'b1010000000000001001000000100000,
31'b0000101000000000001001000100000,
31'b1100000000100000001001000000000,
31'b0000000000000000000100001100000,
31'b0010010000000000000000010001000,
31'b0000001000000000010010000001000,
31'b0010010000000100000000010001000,
31'b0100000100000000000100000000000,
31'b0100000100000010000100000000000,
31'b0100000100000100000100000000000,
31'b0000000010000000100000000000001,
31'b0100000100001000000100000000000,
31'b0101100000000101000000000000000,
31'b0101100000000011000000000000000,
31'b0101100000000001000000000000000,
31'b0000000000000000001000000001001,
31'b1000000000000000100100010000000,
31'b0000000010000000010101000000000,
31'b1100000000000000001001000000000,
31'b0000000000100000000100001100000,
31'b1000010000000000001000001010000,
31'b0000001011000000000000000100001,
31'b1100000000001000001001000000000,
31'b0100000101100000000100000000000,
31'b0100000000000100000000000010100,
31'b0100000000000010000000000010100,
31'b0100000000000000000000000010100,
31'b0101000001000000000000000001100,
31'b0100100000000000000100010000000,
31'b0100100100000000010000000001000,
31'b0100000000001000000000000010100,
31'b0000101000100000000110000000000,
31'b1100000000000000000110000100000,
31'b1100010100000000000000100000000,
31'b1001000000000001100000000000000,
31'b0000100010000000000001000001000,
31'b0110000010000000000000000100100,
31'b0000100010000100000001000001000,
31'b1100100010000000000000000000001,
31'b0100000101000000000100000000000,
31'b0100000101000010000100000000000,
31'b0100000101000100000100000000000,
31'b0100000000100000000000000010100,
31'b1010000100000000010000100000000,
31'b1000010000000000010000010000010,
31'b1010001000000000000010000000010,
31'b0101100001000001000000000000000,
31'b0000101000000000000110000000000,
31'b1001000000000000001010000000010,
31'b0000101000000100000110000000000,
31'b1100000001000000001001000000000,
31'b0000101000001000000110000000000,
31'b0010010000000000010000000010100,
31'b0000001010000000000000000100001,
31'b0001000000000000001000000010001,
31'b1101100000000000000000000000000,
31'b0001001000100000000000000100000,
31'b1101100000000100000000000000000,
31'b0001100000000000000001000001001,
31'b1101100000001000000000000000000,
31'b0010010000000000000010000100100,
31'b0010000100000000000100100000100,
31'b1100000100000001000100000000000,
31'b1101100000010000000000000000000,
31'b0001100100000000100000010000000,
31'b0010000000101000001000000100000,
31'b0000010000000000000000010100001,
31'b0100000000000001001001000000000,
31'b0101001100000000000000001000000,
31'b0010000000100000001000000100000,
31'b1010010000000000000100000010000,
31'b0000000010000000001000000010000,
31'b0001001000000000000000000100000,
31'b0011000000000000000000100001000,
31'b0001001000000100000000000100000,
31'b0001000001010000100000000000000,
31'b0010000001000000000000100010000,
31'b0010000000010000001000000100000,
31'b0010000001000100000000100010000,
31'b0001000001001000100000000000000,
31'b0001001000010000000000000100000,
31'b0010000000001000001000000100000,
31'b0000000000000000100000000011000,
31'b0001000001000000100000000000000,
31'b0001000001000010100000000000000,
31'b0010000000000000001000000100000,
31'b0010000000000010001000000100000,
31'b1101100001000000000000000000000,
31'b0010001000000001000010000000010,
31'b1100000100000000010000000000100,
31'b0010001000100000101000000000000,
31'b0001000000110000100000000000000,
31'b0010000000100000000000100010000,
31'b0001110000000000000000000001010,
31'b1100100000000000000000000011000,
31'b1000000010000000000001000000100,
31'b1001000000000000000000011100000,
31'b1001000000000000010000100000010,
31'b0000000010100000000000100100000,
31'b0001000000100000100000000000000,
31'b0001000000100010100000000000000,
31'b0001000000100100100000000000000,
31'b0001000010000000000000001000110,
31'b0001000000011000100000000000000,
31'b0010000000001000000000100010000,
31'b0011000001000000000000100001000,
31'b0010001000000000101000000000000,
31'b0001000000010000100000000000000,
31'b0010000000000000000000100010000,
31'b0001000000010100100000000000000,
31'b0010000000000100000000100010000,
31'b0001000000001000100000000000000,
31'b0001000000001010100000000000000,
31'b0001000000001100100000000000000,
31'b0000000010000000000000100100000,
31'b0001000000000000100000000000000,
31'b0001000000000010100000000000000,
31'b0001000000000100100000000000000,
31'b0001000000000110100000000000000,
31'b0000000000100000001000000010000,
31'b1000010000000000000100000100000,
31'b1000000100000000000010100000000,
31'b1000010000000100000100000100000,
31'b1000000000000001100000000000001,
31'b1000010000001000000100000100000,
31'b0000001000100000100000100000000,
31'b0100000101000000000000101000000,
31'b1000000001000000000001000000100,
31'b1000010000010000000100000100000,
31'b1000000100010000000010100000000,
31'b0000010000000000000010000010100,
31'b1000000001001000000001000000100,
31'b1000010000000000000000000000111,
31'b0010101000000000010100000000000,
31'b0011001000100000000000000010000,
31'b0000000000000000001000000010000,
31'b0000000000000010001000000010000,
31'b0000000000000100001000000010000,
31'b0000000001010000000000100100000,
31'b0000000000001000001000000010000,
31'b0010000000000000100000000101000,
31'b0000001000000000100000100000000,
31'b0001000001000000001000000001000,
31'b0000000000010000001000000010000,
31'b0000000001000100000000100100000,
31'b0000000001000010000000100100000,
31'b0000000001000000000000100100000,
31'b0001000011000000100000000000000,
31'b0011001000000100000000000010000,
31'b0010000010000000001000000100000,
31'b0011001000000000000000000010000,
31'b1000000000010000000001000000100,
31'b1000010001000000000100000100000,
31'b1000000101000000000010100000000,
31'b0000000100000000001100000000100,
31'b1000000001000001100000000000001,
31'b0110000000000000000010010001000,
31'b0100011000000000010000000001000,
31'b0100000100000000000000101000000,
31'b1000000000000000000001000000100,
31'b1000000000000010000001000000100,
31'b1000000000000100000001000000100,
31'b0000000000100000000000100100000,
31'b1000000000001000000001000000100,
31'b1000000000001010000001000000100,
31'b1000000000001100000001000000100,
31'b0001000000000000000000001000110,
31'b0000000001000000001000000010000,
31'b0000000001000010001000000010000,
31'b0000000001000100001000000010000,
31'b0000000000010000000000100100000,
31'b0001000010010000100000000000000,
31'b0010000010000000000000100010000,
31'b0001000000000010001000000001000,
31'b0001000000000000001000000001000,
31'b0010001000000000000000000001000,
31'b0000000000000100000000100100000,
31'b0000000000000010000000100100000,
31'b0000000000000000000000100100000,
31'b0001000010000000100000000000000,
31'b0001000010000010100000000000000,
31'b0001000010000100100000000000000,
31'b0000000000001000000000100100000,
31'b1101100100000000000000000000000,
31'b0001100000010000100000010000000,
31'b1000000010000000000010100000000,
31'b1100000000001001000100000000000,
31'b0010010000000000001001000010000,
31'b1100000000000101000100000000000,
31'b0010000000000000000100100000100,
31'b1100000000000001000100000000000,
31'b1001001001000000000010000000000,
31'b0001100000000000100000010000000,
31'b1100001000000000000001000000010,
31'b0001100000000100100000010000000,
31'b0101001000000010000000001000000,
31'b0101001000000000000000001000000,
31'b0010000100100000001000000100000,
31'b1100000000010001000100000000000,
31'b0001000000000000000010011000000,
31'b0001001100000000000000000100000,
31'b1100000000000000000000010011000,
31'b0001010000000000000000010001010,
31'b0001000101010000100000000000000,
31'b1101000001000000000000010000000,
31'b0010000100010000001000000100000,
31'b1100000000100001000100000000000,
31'b0001000101001000100000000000000,
31'b0001100000100000100000010000000,
31'b0110000000000000000000000001110,
31'b0000100000000000000001000100010,
31'b0001000101000000100000000000000,
31'b0101001000100000000000001000000,
31'b0010000100000000001000000100000,
31'b0010000100000010001000000100000,
31'b1100000000000100010000000000100,
31'b0010000000000101010000100000000,
31'b1100000000000000010000000000100,
31'b0010000000000001010000100000000,
31'b0001101000000000000000010100000,
31'b1101000000100000000000010000000,
31'b1100000000001000010000000000100,
31'b1010000000000000001010000000000,
31'b1001001000000000000010000000000,
31'b1001001000000010000010000000000,
31'b1100000000010000010000000000100,
31'b0010100000000000001000010100000,
31'b0001000100100000100000000000000,
31'b0101001001000000000000001000000,
31'b0001001000000000000000000010011,
31'b1100011000000000000000000000001,
31'b0001000100011000100000000000000,
31'b1101000000001000000000010000000,
31'b1100000000100000010000000000100,
31'b0010001100000000101000000000000,
31'b0001000100010000100000000000000,
31'b1101000000000000000000010000000,
31'b0001000100010100100000000000000,
31'b1101000000000100000000010000000,
31'b0001000100001000100000000000000,
31'b0101100000000000000010000100000,
31'b0001000100001100100000000000000,
31'b0000100000000001100100000000000,
31'b0001000100000000100000000000000,
31'b0100010000000001000000100000000,
31'b0001000100000100100000000000000,
31'b0101000010000000000100000000001,
31'b1000000000000100000010100000000,
31'b1000010100000000000100000100000,
31'b1000000000000000000010100000000,
31'b1000000000000010000010100000000,
31'b0000000000000101011000000000000,
31'b0100000001000100000000101000000,
31'b0000000000000001011000000000000,
31'b0100000001000000000000101000000,
31'b1000000101000000000001000000100,
31'b0110000000000000100000001001000,
31'b1000000000010000000010100000000,
31'b1000000000100000000101000010000,
31'b0100000000000011000000010000001,
31'b0100000000000001000000010000001,
31'b0000100000000000000000110100000,
31'b0100000001010000000000101000000,
31'b0000000100000000001000000010000,
31'b0000000100000010001000000010000,
31'b1000000000100000000010100000000,
31'b1000000000100010000010100000000,
31'b0000000100001000001000000010000,
31'b0010100000000000000001000010010,
31'b0000001100000000100000100000000,
31'b0101011000000001000000000000000,
31'b0000010001000000000110000000000,
31'b1000010000000000001000100000100,
31'b1000000000110000000010100000000,
31'b1000000000000000000101000010000,
31'b0001000111000000100000000000000,
31'b1100010000000000000100001000000,
31'b0010001000000001000000010000100,
31'b1100001000000000000000110000000,
31'b1000000100010000000001000000100,
31'b0000010000000000000001100010000,
31'b1000000001000000000010100000000,
31'b0000000000000000001100000000100,
31'b0100000000000110000000101000000,
31'b0100000000000100000000101000000,
31'b0100000000000010000000101000000,
31'b0100000000000000000000101000000,
31'b1000000100000000000001000000100,
31'b1000000100000010000001000000100,
31'b1000000100000100000001000000100,
31'b0000000100100000000000100100000,
31'b1010000000000000100010000001000,
31'b0100000001000001000000010000001,
31'b0100100000000000010000000010001,
31'b0100000000010000000000101000000,
31'b0000010000010000000110000000000,
31'b0000010000100000000001100010000,
31'b1000010000000000000000000110100,
31'b0000000100010000000000100100000,
31'b0001000110010000100000000000000,
31'b1101000010000000000000010000000,
31'b0101000000000000110001000000000,
31'b0100000000100000000000101000000,
31'b0000010000000000000110000000000,
31'b0000010000000010000110000000000,
31'b0000010000000100000110000000000,
31'b0000000100000000000000100100000,
31'b0001000110000000100000000000000,
31'b0101000000000100000100000000001,
31'b0101000000000010000100000000001,
31'b0101000000000000000100000000001,
31'b1000000010000000010000000000010,
31'b0001000000100000000000000100000,
31'b1001000000000000000001100000100,
31'b0001000000100100000000000100000,
31'b1001000000000000100000011000000,
31'b0001000000101000000000000100000,
31'b0000000010100000100000100000000,
31'b0001000010000000010001001000000,
31'b1001000101000000000010000000000,
31'b0001000000110000000000000100000,
31'b1100000100000000000001000000010,
31'b0001010100000000000001000010000,
31'b0101000100000010000000001000000,
31'b0101000100000000000000001000000,
31'b0010100010000000010100000000000,
31'b1110100000000000001000000000000,
31'b0001000000000010000000000100000,
31'b0001000000000000000000000100000,
31'b0001000000000110000000000100000,
31'b0001000000000100000000000100000,
31'b0001000000001010000000000100000,
31'b0001000000001000000000000100000,
31'b0000000010000000100000100000000,
31'b0001000000001100000000000100000,
31'b0010000011000000000000000001000,
31'b0001000000010000000000000100000,
31'b0010001000001000001000000100000,
31'b0001000000010100000000000100000,
31'b0001001001000000100000000000000,
31'b0000000000000000001000100001000,
31'b0010001000000000001000000100000,
31'b0011000010000000000000000010000,
31'b1001000100010000000010000000000,
31'b0010000000000001000010000000010,
31'b0010010000000001000000001001000,
31'b0010000000100000101000000000000,
31'b0001100100000000000000010100000,
31'b0010001000100000000000100010000,
31'b0000010000000000100000010000001,
31'b1010000000000001000000000010001,
31'b1001000100000000000010000000000,
31'b1001000100000010000010000000000,
31'b1100100010000000000000100000000,
31'b0010100010000001000000000000100,
31'b0001001000100000100000000000000,
31'b0101000101000000000000001000000,
31'b0001001000100100100000000000000,
31'b1100010100000000000000000000001,
31'b0010000010010000000000000001000,
31'b0001000001000000000000000100000,
31'b0010000000000010101000000000000,
31'b0010000000000000101000000000000,
31'b0001001000010000100000000000000,
31'b0010001000000000000000100010000,
31'b0000000000000000000000000111000,
31'b0010000000001000101000000000000,
31'b0010000010000000000000000001000,
31'b0010000010000010000000000001000,
31'b0010000010000100000000000001000,
31'b0010000000010000101000000000000,
31'b0001001000000000100000000000000,
31'b0001001000000010100000000000000,
31'b0001001000000100100000000000000,
31'b0011000011000000000000000010000,
31'b1000000000000000010000000000010,
31'b1000000000000010010000000000010,
31'b1000000000000100010000000000010,
31'b1000000000000110010000000000010,
31'b1000000000001000010000000000010,
31'b1000000000001010010000000000010,
31'b0000000000100000100000100000000,
31'b0001000000000000010001001000000,
31'b1000000000010000010000000000010,
31'b1000000001000001000000000100001,
31'b1100100001000000000000100000000,
31'b0011000000101000000000000010000,
31'b1000010001000000100100000000000,
31'b0101000110000000000000001000000,
31'b0010100000000000010100000000000,
31'b0011000000100000000000000010000,
31'b0000001000000000001000000010000,
31'b0001000010000000000000000100000,
31'b0000000000001000100000100000000,
31'b0001000010000100000000000100000,
31'b0000000000000100100000100000000,
31'b0001000010001000000000000100000,
31'b0000000000000000100000100000000,
31'b0000000000000010100000100000000,
31'b0010000001000000000000000001000,
31'b0010000001000010000000000001000,
31'b0010000001000100000000000001000,
31'b0011000000001000000000000010000,
31'b0010000001001000000000000001000,
31'b0011000000000100000000000010000,
31'b0000000000010000100000100000000,
31'b0011000000000000000000000010000,
31'b1000000001000000010000000000010,
31'b1000000001000010010000000000010,
31'b1100100000010000000000100000000,
31'b0010100000010001000000000000100,
31'b1000010000010000100100000000000,
31'b1000010000000000010001000000001,
31'b0100010000000000010000000001000,
31'b0100010000000010010000000001000,
31'b0010000000100000000000000001000,
31'b1000000000000001000000000100001,
31'b1100100000000000000000100000000,
31'b0010100000000001000000000000100,
31'b1000010000000000100100000000000,
31'b1000010000000010100100000000000,
31'b1100100000001000000000100000000,
31'b0011000001100000000000000010000,
31'b0010000000010000000000000001000,
31'b0010000000010010000000000001000,
31'b0010000000010100000000000001000,
31'b0010000010000000101000000000000,
31'b0010000000011000000000000001000,
31'b0010001010000000000000100010000,
31'b0000000001000000100000100000000,
31'b0001001000000000001000000001000,
31'b0010000000000000000000000001000,
31'b0010000000000010000000000001000,
31'b0010000000000100000000000001000,
31'b0000001000000000000000100100000,
31'b0010000000001000000000000001000,
31'b0010000000001010000000000001000,
31'b0010000000001100000000000001000,
31'b0011000001000000000000000010000,
31'b1001000001010000000010000000000,
31'b0001000100100000000000000100000,
31'b1100000000010000000001000000010,
31'b0001010000010000000001000010000,
31'b0110100000000000000101000000000,
31'b0101000000010000000000001000000,
31'b0010100000000000101000010000000,
31'b1100001000000001000100000000000,
31'b1001000001000000000010000000000,
31'b0000000000000000000000000001011,
31'b1100000000000000000001000000010,
31'b0001010000000000000001000010000,
31'b0101000000000010000000001000000,
31'b0101000000000000000000001000000,
31'b1100000000001000000001000000010,
31'b1000000000000000000010000011000,
31'b0001000100000010000000000100000,
31'b0001000100000000000000000100000,
31'b0001010000000000000110100000000,
31'b0001000100000100000000000100000,
31'b0101100000000000100010000000000,
31'b0100000000000000000100100000001,
31'b0000100000000001000100000100000,
31'b0101010010000001000000000000000,
31'b1010000000000001000000000100010,
31'b0001000100010000000000000100000,
31'b1100000000100000000001000000010,
31'b0001010000100000000001000010000,
31'b0101000000100010000000001000000,
31'b0101000000100000000000001000000,
31'b0010001100000000001000000100000,
31'b1100000010000000000000110000000,
31'b1001000000010000000010000000000,
31'b1010000000100000010000000000001,
31'b1100001000000000010000000000100,
31'b0010001000000001010000100000000,
31'b0001100000000000000000010100000,
31'b0101000001010000000000001000000,
31'b0001100000000100000000010100000,
31'b1100010000010000000000000000001,
31'b1001000000000000000010000000000,
31'b1001000000000010000010000000000,
31'b1001000000000100000010000000000,
31'b1100010000001000000000000000001,
31'b0000010000000000000001000001000,
31'b0101000001000000000000001000000,
31'b0001000000000000000000000010011,
31'b1100010000000000000000000000001,
31'b1010000000000010010000000000001,
31'b1010000000000000010000000000001,
31'b0110000000000000010001000001000,
31'b0010000100000000101000000000000,
31'b0001100000100000000000010100000,
31'b1101001000000000000000010000000,
31'b0000100000000000100001000000010,
31'b0010000100001000101000000000000,
31'b1001000000100000000010000000000,
31'b1010000000010000010000000000001,
31'b1110000000000000001000010000000,
31'b0010000100010000101000000000000,
31'b0001001100000000100000000000000,
31'b0101000001100000000000001000000,
31'b0001001100000100100000000000000,
31'b1100010000100000000000000000001,
31'b1000000100000000010000000000010,
31'b1010000000000000000010000101000,
31'b1000001000000000000010100000000,
31'b1000001000000010000010100000000,
31'b1000000100001000010000000000010,
31'b0101000010010000000000001000000,
31'b0000001000000001011000000000000,
31'b0101010000100001000000000000000,
31'b1001000011000000000010000000000,
31'b0011000000000001010000000000000,
31'b1100000010000000000001000000010,
31'b0011000000000101010000000000000,
31'b0101000010000010000000001000000,
31'b0101000010000000000000001000000,
31'b0010100100000000010100000000000,
31'b1100000000100000000000110000000,
31'b0000000000000001000010000000001,
31'b0001000110000000000000000100000,
31'b0000000100001000100000100000000,
31'b0101010000001001000000000000000,
31'b0000000100000100100000100000000,
31'b0101010000000101000000000000000,
31'b0000000100000000100000100000000,
31'b0101010000000001000000000000000,
31'b0010000101000000000000000001000,
31'b0011000000100001010000000000000,
31'b0010000101000100000000000001000,
31'b1100000000001000000000110000000,
31'b0010000101001000000000000001000,
31'b1100000000000100000000110000000,
31'b0010000000000001000000010000100,
31'b1100000000000000000000110000000,
31'b1001000010010000000010000000000,
31'b0100010000001000000100010000000,
31'b1001100000000000000000000000110,
31'b0000100000000000100000110000000,
31'b0110000000000000000000001101000,
31'b0100010000000000000100010000000,
31'b0100010100000000010000000001000,
31'b0100001000000000000000101000000,
31'b1001000010000000000010000000000,
31'b1001000010000010000010000000000,
31'b1100100100000000000000100000000,
31'b0010100100000001000000000000100,
31'b0011000000000000000100000000100,
31'b0101000011000000000000001000000,
31'b0011000000000100000100000000100,
31'b1100010010000000000000000000001,
31'b0010000100010000000000000001000,
31'b1010000010000000010000000000001,
31'b0010000100010100000000000001000,
31'b0010000110000000101000000000000,
31'b0010000100011000000000000001000,
31'b1100000000000001000000001000001,
31'b0000000101000000100000100000000,
31'b0101010001000001000000000000000,
31'b0010000100000000000000000001000,
31'b0010000100000010000000000001000,
31'b0010000100000100000000000001000,
31'b0010000000000000010100010000000,
31'b0010000100001000000000000001000,
31'b0010100000000000010000000010100,
31'b0010000100001100000000000001000,
31'b1100000001000000000000110000000,
31'b0100000000000000011000000100000,
31'b0000100000000000000000000010010,
31'b0100100001000000000000001000001,
31'b0000100000000100000000000010010,
31'b0100100000000000000011000001000,
31'b0010000000000000000010000100100,
31'b1001000000000000100100100000000,
31'b1000100000000000000010000000001,
31'b0100100000000001000000110000000,
31'b0000100000010000000000000010010,
31'b0000000000000010000000010100001,
31'b0000000000000000000000010100001,
31'b0101000000000000010000100001000,
31'b1010000000000100000100000010000,
31'b1010000000000010000100000010000,
31'b1010000000000000000100000010000,
31'b0001000000000000010100000000010,
31'b0001011000000000000000000100000,
31'b0011010000000000000000100001000,
31'b0001011000000100000000000100000,
31'b0001010001010000100000000000000,
31'b0010010001000000000000100010000,
31'b1010000000000000000011100000000,
31'b1000100000100000000010000000001,
31'b0001010001001000100000000000000,
31'b0001011000010000000000000100000,
31'b1010000000000001000000010001000,
31'b0000010000000000100000000011000,
31'b0001010001000000100000000000000,
31'b0100000101000001000000100000000,
31'b1000000000000000100000001000001,
31'b1010000000100000000100000010000,
31'b0100100000000100000000001000001,
31'b0000100001000000000000000010010,
31'b0100100000000000000000001000001,
31'b0100100000000010000000001000001,
31'b0001100000000100000000000001010,
31'b0010010000100000000000100010000,
31'b0001100000000000000000000001010,
31'b1000100001000000000010000000001,
31'b1011000000000000000100000001000,
31'b0100000000000100010000100010000,
31'b0100100000010000000000001000001,
31'b0100000000000000010000100010000,
31'b0001010000100000100000000000000,
31'b0100001000000000111000000000000,
31'b0001100000010000000000000001010,
31'b1100001100000000000000000000001,
31'b0001010000011000100000000000000,
31'b0010101000000000000000001000100,
31'b1000000100000000000010010000001,
31'b1000001000000000000000001100001,
31'b0001010000010000100000000000000,
31'b0010010000000000000000100010000,
31'b0001100000100000000000000001010,
31'b0010010000000100000000100010000,
31'b0001010000001000100000000000000,
31'b0100000100001001000000100000000,
31'b0101100000000000000100100000000,
31'b0100000000000000100010000000001,
31'b0001010000000000100000000000000,
31'b0100000100000001000000100000000,
31'b0001010000000100100000000000000,
31'b0100000100000101000000100000000,
31'b1000000000000010000100000100000,
31'b1000000000000000000100000100000,
31'b1000010100000000000010100000000,
31'b1000000000000100000100000100000,
31'b1000010000000001100000000000001,
31'b1000000000001000000100000100000,
31'b0100001001000000010000000001000,
31'b1000100010000000000010000000001,
31'b1000010001000000000001000000100,
31'b1000000000010000000100000100000,
31'b0000000100000000001001000100000,
31'b0000000000000000000010000010100,
31'b1000001001000000100100000000000,
31'b1000000000000000000000000000111,
31'b0110000000000000011000000010000,
31'b0010100000000000000000000100010,
31'b0000010000000000001000000010000,
31'b1000000000100000000100000100000,
31'b0000010000000100001000000010000,
31'b1000000001000000001011000000000,
31'b0000010000001000001000000010000,
31'b1000000000101000000100000100000,
31'b0100000000000000001001001000000,
31'b0101001100000001000000000000000,
31'b0000010000010000001000000010000,
31'b1000000100000000001000100000100,
31'b0000010001000010000000100100000,
31'b0000010001000000000000100100000,
31'b0001010011000000100000000000000,
31'b1100000100000000000100001000000,
31'b1110001000000000000000000000010,
31'b0011011000000000000000000010000,
31'b1000010000010000000001000000100,
31'b1000000001000000000100000100000,
31'b0100100010000000000000001000001,
31'b1000000001000100000100000100000,
31'b1000001000010000100100000000000,
31'b1000001000000000010001000000001,
31'b0100001000000000010000000001000,
31'b0100010100000000000000101000000,
31'b1000010000000000000001000000100,
31'b1000010000000010000001000000100,
31'b1000010000000100000001000000100,
31'b0000010000100000000000100100000,
31'b1000001000000000100100000000000,
31'b1000001000000010100100000000000,
31'b1100000000000000000000001010100,
31'b0010100001000000000000000100010,
31'b0000010001000000001000000010000,
31'b1000000001100000000100000100000,
31'b1000000100000000000000000110100,
31'b1000000000000000001011000000000,
31'b0001010010010000100000000000000,
31'b0010010010000000000000100010000,
31'b0100001000100000010000000001000,
31'b0001010000000000001000000001000,
31'b0000000100000000000110000000000,
31'b0000010000000100000000100100000,
31'b0000010000000010000000100100000,
31'b0000010000000000000000100100000,
31'b0001010010000000100000000000000,
31'b0100100000000000100100000100000,
31'b0001100000000011000010000000000,
31'b0001100000000001000010000000000,
31'b0110100000000000100000000000100,
31'b0000100100000000000000000010010,
31'b1100000000000000100000000100001,
31'b0001001000010000000001000010000,
31'b0010000000000000001001000010000,
31'b0010000100000000000010000100100,
31'b0010010000000000000100100000100,
31'b1100010000000001000100000000000,
31'b0000001001001000000001000001000,
31'b0001110000000000100000010000000,
31'b0000001000000000000010001000001,
31'b0001001000000000000001000010000,
31'b0000001001000000000001000001000,
31'b0101011000000000000000001000000,
31'b0000100010000000010010000001000,
31'b1100001001000000000000000000001,
31'b0001010000000000000010011000000,
31'b0001011100000000000000000100000,
31'b1000000001000000000010010000001,
31'b0001000000000000000000010001010,
31'b0000000001000000000000010010010,
31'b0100000001010001000000100000000,
31'b0100000000000010000000011000001,
31'b0100000000000000000000011000001,
31'b0000000011000000000110000000000,
31'b1010000000000001010100000000000,
31'b0000101000000000010101000000000,
31'b0001001000100000000001000010000,
31'b0000000000000000011000001000000,
31'b0100000001000001000000100000000,
31'b0000100001000000000000000100001,
31'b0100000001000101000000100000000,
31'b0000001000011000000001000001000,
31'b0000000010000000000001100010000,
31'b1100010000000000010000000000100,
31'b0011000000000000001001000001000,
31'b0000001000010000000001000001000,
31'b0100001010000000000100010000000,
31'b0001100100000000000000000001010,
31'b1100001000010000000000000000001,
31'b0000001000001000000001000001000,
31'b0100001000000000000010000010010,
31'b0000100000101000000000000100001,
31'b1100001000001000000000000000001,
31'b0000001000000000000001000001000,
31'b0100000000100001000000100000000,
31'b0000100000100000000000000100001,
31'b1100001000000000000000000000001,
31'b0000000010010000000110000000000,
31'b0100000000011001000000100000000,
31'b1000000000000000000010010000001,
31'b1001001000000000001000000000100,
31'b0000000000000000000000010010010,
31'b0100000000010001000000100000000,
31'b0000100000010000000000000100001,
31'b0100000001000000000000011000001,
31'b0000000010000000000110000000000,
31'b0100000000001001000000100000000,
31'b0000100000001000000000000100001,
31'b0100000100000000100010000000001,
31'b1010000000000000000000000000100,
31'b0100000000000001000000100000000,
31'b0000100000000000000000000100001,
31'b0100000000000101000000100000000,
31'b1000010000000100000010100000000,
31'b1000000100000000000100000100000,
31'b1000010000000000000010100000000,
31'b1000010000000010000010100000000,
31'b0011000000000001000000000000101,
31'b1101000000000000000000100000001,
31'b0001000000000000000001100001000,
31'b0101001000100001000000000000000,
31'b0000000001100000000110000000000,
31'b1000000100010000000100000100000,
31'b0000000000000000001001000100000,
31'b0000000100000000000010000010100,
31'b0000101000000000000100001100000,
31'b1100000000100000000100001000000,
31'b0000100000000000010010000001000,
31'b0010100100000000000000000100010,
31'b0000010100000000001000000010000,
31'b1000000100100000000100000100000,
31'b1000010000100000000010100000000,
31'b0110100000000000000000001000010,
31'b0000010100001000001000000010000,
31'b1100000000010000000100001000000,
31'b0101001000000011000000000000000,
31'b0101001000000001000000000000000,
31'b0000000001000000000110000000000,
31'b1000000000000000001000100000100,
31'b0000000001000100000110000000000,
31'b1000010000000000000101000010000,
31'b0000000010000000011000001000000,
31'b1100000000000000000100001000000,
31'b0000100011000000000000000100001,
31'b1100000000000100000100001000000,
31'b0000000000110000000110000000000,
31'b0000000000000000000001100010000,
31'b1000010001000000000010100000000,
31'b0000010000000000001100000000100,
31'b0100001000000010000100010000000,
31'b0100001000000000000100010000000,
31'b0100010000000010000000101000000,
31'b0100010000000000000000101000000,
31'b0000000000100000000110000000000,
31'b0000000000100010000110000000000,
31'b0000000001000000001001000100000,
31'b0000010100100000000000100100000,
31'b0000001010000000000001000001000,
31'b0100001000010000000100010000000,
31'b0000100010100000000000000100001,
31'b1100001010000000000000000000001,
31'b0000000000010000000110000000000,
31'b0000000000100000000001100010000,
31'b1000000000000000000000000110100,
31'b1000000100000000001011000000000,
31'b0000000010000000000000010010010,
31'b0100001000100000000100010000000,
31'b1010100000000000000010000000010,
31'b0101001001000001000000000000000,
31'b0000000000000000000110000000000,
31'b0000000000000010000110000000000,
31'b0000000000000100000110000000000,
31'b0000010100000000000000100100000,
31'b0000000000001000000110000000000,
31'b0100000010000001000000100000000,
31'b0000100010000000000000000100001,
31'b0101010000000000000100000000001,
31'b1001000000000000001100000010000,
31'b0001010000100000000000000100000,
31'b0010000100000000100001100000000,
31'b0001010000100100000000000100000,
31'b0010000100000000000000011000100,
31'b0011000000000001000000001010000,
31'b0000000001000000100000010000001,
31'b1000101000000000000010000000001,
31'b0010000001000000100010000000100,
31'b0001010000110000000000000100000,
31'b0000000100000000000010001000001,
31'b0001000100000000000001000010000,
31'b0000000101000000000001000001000,
31'b0101010100000000000000001000000,
31'b0000000101000100000001000001000,
31'b1100000101000000000000000000001,
31'b0100100010000000000100000000000,
31'b0001010000000000000000000100000,
31'b0100100010000100000100000000000,
31'b0001010000000100000000000100000,
31'b0100100010001000000100000000000,
31'b0001010000001000000000000100000,
31'b0100000000000000000010000100001,
31'b0101000110000001000000000000000,
31'b0110000000000000000000010100100,
31'b0001010000010000000000000100000,
31'b1100100000000000000000010000001,
31'b0001010000010100000000000100000,
31'b0001011001000000100000000000000,
31'b0001000000000001010001000000000,
31'b1110000010000000000000000000010,
31'b0011010010000000000000000010000,
31'b0010000000010000100010000000100,
31'b0010100000100000000000001000100,
31'b0010000000000001000000001001000,
31'b1000000000100000000000001100001,
31'b0000000100010000000001000001000,
31'b1000000010000000010001000000001,
31'b0000000000000000100000010000001,
31'b1000000000000000001100000001000,
31'b0010000000000000100010000000100,
31'b0100000100000000000010000010010,
31'b0010000000010001000000001001000,
31'b1100000100001000000000000000001,
31'b0000000100000000000001000001000,
31'b0100000000000000111000000000000,
31'b0000000100000100000001000001000,
31'b1100000100000000000000000000001,
31'b0100100011000000000100000000000,
31'b0010100000000000000000001000100,
31'b1000000000000010000000001100001,
31'b1000000000000000000000001100001,
31'b0001011000010000100000000000000,
31'b0010100000001000000000001000100,
31'b0000010000000000000000000111000,
31'b1000000000100000001100000001000,
31'b0010010010000000000000000001000,
31'b0010100000010000000000001000100,
31'b0010010010000100000000000001000,
31'b1100000000000000001000100000010,
31'b0001011000000000100000000000000,
31'b0100001100000001000000100000000,
31'b0001100000000000000001010010000,
31'b1100000100100000000000000000001,
31'b1000010000000000010000000000010,
31'b1000001000000000000100000100000,
31'b1010000000000000000100100001000,
31'b1000001000000100000100000100000,
31'b1000010000001000010000000000010,
31'b1000001000001000000100000100000,
31'b0100000001000000010000000001000,
31'b0101000100100001000000000000000,
31'b1000010000010000010000000000010,
31'b1000001000010000000100000100000,
31'b0001000000000011000000001100000,
31'b0001000000000001000000001100000,
31'b1000000001000000100100000000000,
31'b1000001000000000000000000000111,
31'b1110000000100000000000000000010,
31'b0011010000100000000000000010000,
31'b0100100000000000000100000000000,
31'b0100100000000010000100000000000,
31'b0100100000000100000100000000000,
31'b0101000100001001000000000000000,
31'b0100100000001000000100000000000,
31'b0101000100000101000000000000000,
31'b0000010000000000100000100000000,
31'b0101000100000001000000000000000,
31'b0100100000010000000100000000000,
31'b0111000000000000000001001000000,
31'b1110000000001000000000000000010,
31'b0011010000001000000000000010000,
31'b1110000000000100000000000000010,
31'b0011010000000100000000000010000,
31'b1110000000000000000000000000010,
31'b0011010000000000000000000010000,
31'b1000010001000000010000000000010,
31'b1000001001000000000100000100000,
31'b0100000000001000010000000001000,
31'b0100100100000000000000000010100,
31'b1000000000010000100100000000000,
31'b1000000000000000010001000000001,
31'b0100000000000000010000000001000,
31'b0100000000000010010000000001000,
31'b1000000000001000100100000000000,
31'b1000010000000001000000000100001,
31'b1100110000000000000000100000000,
31'b0010110000000001000000000000100,
31'b1000000000000000100100000000000,
31'b1000000000000010100100000000000,
31'b1000000000000100100100000000000,
31'b1100000110000000000000000000001,
31'b0100100001000000000100000000000,
31'b0101000000000000000000010001100,
31'b0100100001000100000100000000000,
31'b1000001000000000001011000000000,
31'b1010100000000000010000100000000,
31'b1000100000000000000110001000000,
31'b0100000000100000010000000001000,
31'b0101000101000001000000000000000,
31'b0010010000000000000000000001000,
31'b0010010000000010000000000001000,
31'b0010010000000100000000000001000,
31'b0010000000000000000010001000010,
31'b1000000000100000100100000000000,
31'b1010000000000000000000001010001,
31'b1110000001000000000000000000010,
31'b0011010001000000000000000010000,
31'b0010000000001000000000011000100,
31'b0001010100100000000000000100000,
31'b0010000000000000100001100000000,
31'b0001000000010000000001000010000,
31'b0010000000000000000000011000100,
31'b0101010000010000000000001000000,
31'b0010000000001000100001100000000,
31'b1100000001010000000000000000001,
31'b0000000001001000000001000001000,
31'b0001000000000100000001000010000,
31'b0000000000000000000010001000001,
31'b0001000000000000000001000010000,
31'b0000000001000000000001000001000,
31'b0101010000000000000000001000000,
31'b0000000001000100000001000001000,
31'b1100000001000000000000000000001,
31'b0100100110000000000100000000000,
31'b0001010100000000000000000100000,
31'b0001000000000000000110100000000,
31'b0000100000000000100000000000001,
31'b1010000000000000010001000000010,
31'b0101000010000101000000000000000,
31'b0101000010000011000000000000000,
31'b0101000010000001000000000000000,
31'b0000100010000000001000000001001,
31'b0001010100010000000000000100000,
31'b0000100000000000010101000000000,
31'b0001000000100000000001000010000,
31'b0000001000000000011000001000000,
31'b0101010000100000000000001000000,
31'b0000101001000000000000000100001,
31'b1100000001100000000000000000001,
31'b0000000000011000000001000001000,
31'b0100000010001000000100010000000,
31'b0010000100000001000000001001000,
31'b1100000000011000000000000000001,
31'b0000000000010000000001000001000,
31'b0100000010000000000100010000000,
31'b0000000100000000100000010000001,
31'b1100000000010000000000000000001,
31'b0000000000001000000001000001000,
31'b0100000000000000000010000010010,
31'b0000000001000000000010001000001,
31'b1100000000001000000000000000001,
31'b0000000000000000000001000001000,
31'b0000000000000010000001000001000,
31'b0000000000000100000001000001000,
31'b1100000000000000000000000000001,
31'b0100000010000001000000000011000,
31'b1010010000000000010000000000001,
31'b1001000000000010001000000000100,
31'b1001000000000000001000000000100,
31'b0000001000000000000000010010010,
31'b0100001000010001000000100000000,
31'b0000110000000000100001000000010,
31'b1100000000110000000000000000001,
31'b0000001010000000000110000000000,
31'b0100001000001001000000100000000,
31'b0000101000001000000000000100001,
31'b1100000000101000000000000000001,
31'b0000000000100000000001000001000,
31'b0100001000000001000000100000000,
31'b0000101000000000000000000100001,
31'b1100000000100000000000000000001,
31'b1000010100000000010000000000010,
31'b1010000000000000010000110000000,
31'b1010000000000000000000001100010,
31'b0101000000101001000000000000000,
31'b0101100000000000000000000001100,
31'b0100000001000000000100010000000,
31'b0101000000100011000000000000000,
31'b0101000000100001000000000000000,
31'b0000100000100000001000000001001,
31'b0011010000000001010000000000000,
31'b0000001000000000001001000100000,
31'b0001000010000000000001000010000,
31'b0000100000000000000100001100000,
31'b0101010010000000000000001000000,
31'b0000101000000000010010000001000,
31'b1100000011000000000000000000001,
31'b0100100100000000000100000000000,
31'b0101000000001101000000000000000,
31'b0101000000001011000000000000000,
31'b0101000000001001000000000000000,
31'b0101000000000111000000000000000,
31'b0101000000000101000000000000000,
31'b0101000000000011000000000000000,
31'b0101000000000001000000000000000,
31'b0000100000000000001000000001001,
31'b1000100000000000100100010000000,
31'b0000100010000000010101000000000,
31'b1100100000000000001001000000000,
31'b0000100000100000000100001100000,
31'b1100001000000000000100001000000,
31'b1110000100000000000000000000010,
31'b1000000000000000100000000010100,
31'b0100000000100001000000000011000,
31'b0100000000001000000100010000000,
31'b0100100000000010000000000010100,
31'b0100100000000000000000000010100,
31'b0100000000000010000100010000000,
31'b0100000000000000000100010000000,
31'b0100000100000000010000000001000,
31'b0000000000000000101001000000000,
31'b0000001000100000000110000000000,
31'b0100000010000000000010000010010,
31'b0000001001000000001001000100000,
31'b1100000010001000000000000000001,
31'b0000000010000000000001000001000,
31'b0100000000010000000100010000000,
31'b0000000010000100000001000001000,
31'b1100000010000000000000000000001,
31'b0100000000000001000000000011000,
31'b0100000000101000000100010000000,
31'b1001000000000001000010001000000,
31'b1001000010000000001000000000100,
31'b0100000000100010000100010000000,
31'b0100000000100000000100010000000,
31'b0101000001000011000000000000000,
31'b0101000001000001000000000000000,
31'b0000001000000000000110000000000,
31'b0000001000000010000110000000000,
31'b0000001000000100000110000000000,
31'b0010010000000000010100010000000,
31'b0000001000001000000110000000000,
31'b0100001010000001000000100000000,
31'b0000101010000000000000000100001,
31'b1100000010100000000000000000001,
31'b1110000000000000000000000000000,
31'b0000000000000001000000100000100,
31'b1110000000000100000000000000000,
31'b0010000000000000000001000001001,
31'b1110000000001000000000000000000,
31'b0010000001000000000010001000000,
31'b1110000000001100000000000000000,
31'b0010000001000100000010001000000,
31'b1110000000010000000000000000000,
31'b0010000100000000100000010000000,
31'b1110000000010100000000000000000,
31'b0010000100000100100000010000000,
31'b1110000000011000000000000000000,
31'b0010000100001000100000010000000,
31'b1000010000100000010000000000000,
31'b1101001000000000001000000000000,
31'b1110000000100000000000000000000,
31'b0010101000000000000000000100000,
31'b0000100000000000000000100001000,
31'b1000001000000000000000000000101,
31'b1110000000101000000000000000000,
31'b0010101000001000000000000100000,
31'b1000010000010000010000000000000,
31'b1000010000010010010000000000000,
31'b1110000000110000000000000000000,
31'b0010101000010000000000000100000,
31'b1000010000001000010000000000000,
31'b1000010000001010010000000000000,
31'b1000010000000100010000000000000,
31'b1010001000000000000010010000000,
31'b1000010000000000010000000000000,
31'b1000010000000010010000000000000,
31'b1110000001000000000000000000000,
31'b0010000000001000000010001000000,
31'b1110000001000100000000000000000,
31'b0010000001000000000001000001001,
31'b0000000000000000010100100000000,
31'b0010000000000000000010001000000,
31'b0010010000000000000000000001010,
31'b0010000000000100000010001000000,
31'b1110000001010000000000000000000,
31'b0010000101000000100000010000000,
31'b0001001000000000001010001000000,
31'b0000000100000001000011000000000,
31'b0010100000100000100000000000000,
31'b0010000000010000000010001000000,
31'b1100000000000000100000100001000,
31'b0010000000010100000010001000000,
31'b1110000001100000000000000000000,
31'b0010101001000000000000000100000,
31'b1000000000000000100100000000010,
31'b1000001001000000000000000000101,
31'b0010100000010000100000000000000,
31'b0010000000100000000010001000000,
31'b1000010001010000010000000000000,
31'b0101000000000000001000011000000,
31'b0100000000000000010000000001010,
31'b0110000100000000000010000100000,
31'b1000010001001000010000000000000,
31'b1000010000000001000100000000100,
31'b0010100000000000100000000000000,
31'b0010100000000010100000000000000,
31'b1000010001000000010000000000000,
31'b1000010001000010010000000000000,
31'b1110000010000000000000000000000,
31'b0010000000000000011100000000000,
31'b1110000010000100000000000000000,
31'b0010000010000000000001000001001,
31'b1000000000000001010000001000000,
31'b1100000001000000001000100000000,
31'b1100000000010000000000000110000,
31'b0001010000010000000000000100010,
31'b1110000010010000000000000000000,
31'b0010000110000000100000010000000,
31'b1100000000001000000000000110000,
31'b0001010000001000000000000100010,
31'b1100000000000100000000000110000,
31'b0001010000000100000000000100010,
31'b1100000000000000000000000110000,
31'b0001010000000000000000000100010,
31'b1110000010100000000000000000000,
31'b0010101010000000000000000100000,
31'b1000000100000000000000001010000,
31'b1000001010000000000000000000101,
31'b1100010100000000000001000000000,
31'b0001100000000000100000000101000,
31'b1000010010010000010000000000000,
31'b0000101000010000000000000010000,
31'b0001101001000000000000000001000,
31'b0000100000000000101000100000000,
31'b1000010010001000010000000000000,
31'b0000101000001000000000000010000,
31'b1010000000000001000001000010000,
31'b0000101000000100000000000010000,
31'b1000010010000000010000000000000,
31'b0000101000000000000000000010000,
31'b1110000011000000000000000000000,
31'b1000000000000000000100001000100,
31'b0001011000000000100000000000010,
31'b1100001000000000100000000010000,
31'b0010000000000001001000000000100,
31'b1100000000000000001000100000000,
31'b0010010010000000000000000001010,
31'b1100000000000100001000100000000,
31'b0001101000100000000000000001000,
31'b1101000000000000000000000101000,
31'b0001000000000000000001000100001,
31'b0001001000000001000000000000100,
31'b0010100010100000100000000000000,
31'b1100000000010000001000100000000,
31'b1100000001000000000000000110000,
31'b0010100000000000000000001000110,
31'b0001101000010000000000000001000,
31'b1100000100000000000000000000011,
31'b0000100000000000100000000110000,
31'b0100000100001000000010000010000,
31'b0010100010010000100000000000000,
31'b1100000000100000001000100000000,
31'b0100000100000010000010000010000,
31'b0100000100000000000010000010000,
31'b0001101000000000000000000001000,
31'b1001000000000000000000100000101,
31'b0001101000000100000000000001000,
31'b0011100000000000000000100100000,
31'b0010100010000000100000000000000,
31'b0010100010000010100000000000000,
31'b1000010011000000010000000000000,
31'b0010010000000001000010000000000,
31'b1110000100000000000000000000000,
31'b0010000000010000100000010000000,
31'b1110000100000100000000000000000,
31'b0010000100000000000001000001001,
31'b1110000100001000000000000000000,
31'b0010000101000000000010001000000,
31'b0001100000000000000100100000100,
31'b0000000001000000000000110001000,
31'b1000010000000001000000000010000,
31'b0010000000000000100000010000000,
31'b1010000010000000010001000000000,
31'b0010000000000100100000010000000,
31'b1010000000100000000000001100000,
31'b0010000000001000100000010000000,
31'b1100000000000001000001001000000,
31'b0010000000001100100000010000000,
31'b1110000100100000000000000000000,
31'b0010101100000000000000000100000,
31'b1000000010000000000000001010000,
31'b1000001100000000000000000000101,
31'b1100010010000000000001000000000,
31'b0001000010000000000001000010010,
31'b1000010100010000010000000000000,
31'b0000010010000000000000000001001,
31'b1010000000001000000000001100000,
31'b0010000000100000100000010000000,
31'b1000010100001000010000000000000,
31'b0101000000000000101010000000000,
31'b1010000000000000000000001100000,
31'b1010000000000010000000001100000,
31'b1000010100000000010000000000000,
31'b1000010100000010010000000000000,
31'b1110000101000000000000000000000,
31'b0010000100001000000010001000000,
31'b0000001010010000000000010010000,
31'b0000000000010001000011000000000,
31'b0010001000000000000000010100000,
31'b0010000100000000000010001000000,
31'b0000001000000000000110000000010,
31'b0000000000000000000000110001000,
31'b1010101000000000000010000000000,
31'b0010000001000000100000010000000,
31'b0000001010000000000000010010000,
31'b0000000000000001000011000000000,
31'b0010100100100000100000000000000,
31'b0010000100010000000010001000000,
31'b0100000010000000000101100000000,
31'b0000000000010000000000110001000,
31'b0001010010000000000000000010001,
31'b1100000010000000000000000000011,
31'b0000000010000000000001000001010,
31'b0100000010001000000010000010000,
31'b0010100100010000100000000000000,
31'b1110100000000000000000010000000,
31'b0100001000000001000001010000000,
31'b0100000010000000000010000010000,
31'b0110000000000010000010000100000,
31'b0110000000000000000010000100000,
31'b0100001000000000000010100001000,
31'b0100000000000000000100010000010,
31'b0010100100000000100000000000000,
31'b0110000000001000000010000100000,
31'b1001000000000000101000001000000,
31'b0100000010010000000010000010000,
31'b1110000110000000000000000000000,
31'b0010000100000000011100000000000,
31'b1000000000100000000000001010000,
31'b1010000000000000100100000000001,
31'b1100010000100000000001000000000,
31'b0001001000010000000000010001000,
31'b1010010000000001000000000100000,
31'b0000010000100000000000000001001,
31'b1010000000000100010001000000000,
31'b0010000010000000100000010000000,
31'b1010000000000000010001000000000,
31'b1010000000000010010001000000000,
31'b0001001000000010000000010001000,
31'b0001001000000000000000010001000,
31'b1100000100000000000000000110000,
31'b0001010100000000000000000100010,
31'b1000000000000100000000001010000,
31'b1100000001000000000000000000011,
31'b1000000000000000000000001010000,
31'b1000000000000010000000001010000,
31'b1100010000000000000001000000000,
31'b0001000000000000000001000010010,
31'b1000000000001000000000001010000,
31'b0000010000000000000000000001001,
31'b1100000000000001010000000100000,
31'b0010000010100000100000010000000,
31'b1000000000010000000000001010000,
31'b1000100000000000010000100000001,
31'b1100010000010000000001000000000,
31'b0001001000100000000000010001000,
31'b1000010110000000010000000000000,
31'b0000101100000000000000000010000,
31'b0001010000100000000000000010001,
31'b1100000000100000000000000000011,
31'b0000001000010000000000010010000,
31'b0100001000000001000000100000010,
31'b0010001010000000000000010100000,
31'b1100000100000000001000100000000,
31'b0100000000100010000010000010000,
31'b0100000000100000000010000010000,
31'b0000110000000000100001000000000,
31'b0010010000000000010010000010000,
31'b0000001000000000000000010010000,
31'b0000001000000010000000010010000,
31'b0000101000000000000100000000100,
31'b1001000000000000001000000000110,
31'b0100000000000000000101100000000,
31'b0100000000110000000010000010000,
31'b0001010000000000000000000010001,
31'b1100000000000000000000000000011,
31'b0000000000000000000001000001010,
31'b0100000000001000000010000010000,
31'b1100010001000000000001000000000,
31'b1001000000000000000000001001000,
31'b0100000000000010000010000010000,
31'b0100000000000000000010000010000,
31'b0001101100000000000000000001000,
31'b1100000000010000000000000000011,
31'b0000001000100000000000010010000,
31'b0100000010000000000100010000010,
31'b0010100110000000100000000000000,
31'b1100000000000000000100000100100,
31'b0100000000100000000101100000000,
31'b0100000000010000000010000010000,
31'b1110001000000000000000000000000,
31'b0010100000100000000000000100000,
31'b1110001000000100000000000000000,
31'b1000000000100000000000000000101,
31'b1110001000001000000000000000000,
31'b0010100000101000000000000100000,
31'b0001000100000000101000010000000,
31'b1101000000010000001000000000000,
31'b1110001000010000000000000000000,
31'b0010100000110000000000000100000,
31'b0001000010001000010100000000000,
31'b1101000000001000001000000000000,
31'b0001000010000100010100000000000,
31'b1101000000000100001000000000000,
31'b0001000010000000010100000000000,
31'b1101000000000000001000000000000,
31'b0100000000000000000001000001100,
31'b0010100000000000000000000100000,
31'b1000000000000010000000000000101,
31'b1000000000000000000000000000101,
31'b0110000100000000100010000000000,
31'b0010100000001000000000000100000,
31'b1000011000010000010000000000000,
31'b1000000000001000000000000000101,
31'b0110000001000000000000011000000,
31'b0010100000010000000000000100000,
31'b1000011000001000010000000000000,
31'b1000000000010000000000000000101,
31'b1010000000000010000010010000000,
31'b1010000000000000000010010000000,
31'b1000011000000000010000000000000,
31'b0000100010000000000000000010000,
31'b1110001001000000000000000000000,
31'b0010100001100000000000000100000,
31'b0001010010000000100000000000010,
31'b1100000010000000100000000010000,
31'b0010000100000000000000010100000,
31'b0010001000000000000010001000000,
31'b0000010000000000010000011000000,
31'b0010001000000100000010001000000,
31'b1100000000000000001000000011000,
31'b0001010000000000001000000001010,
31'b0001000000000000001010001000000,
31'b0001000010000001000000000000100,
31'b0010101000100000100000000000000,
31'b1110000000000000100000000100000,
31'b0001000011000000010100000000000,
31'b1101000001000000001000000000000,
31'b0110000000010000000000011000000,
31'b0010100001000000000000000100000,
31'b1000001000000000100100000000010,
31'b1000000001000000000000000000101,
31'b0010101000010000100000000000000,
31'b0010100001001000000000000100000,
31'b1000010000000000000001000000110,
31'b1000000001001000000000000000101,
31'b0110000000000000000000011000000,
31'b0110000000000010000000011000000,
31'b0110000000000100000000011000000,
31'b1000000001010000000000000000101,
31'b0010101000000000100000000000000,
31'b1010000001000000000010010000000,
31'b1000011001000000010000000000000,
31'b1000000000000001100001000000000,
31'b1110001010000000000000000000000,
31'b0010100010100000000000000100000,
31'b0001010001000000100000000000010,
31'b1100000001000000100000000010000,
31'b1101000000000000100000000001000,
31'b0001000100010000000000010001000,
31'b0001000000010000010100000000000,
31'b0001000000000000100001000000001,
31'b0001100001100000000000000001000,
31'b0000100100000001010000000000000,
31'b0001000000001000010100000000000,
31'b0001000001000001000000000000100,
31'b0001000000000100010100000000000,
31'b0001000100000000000000010001000,
31'b0001000000000000010100000000000,
31'b0000100000100000000000000010000,
31'b0111010000000000000100000000000,
31'b0010100010000000000000000100000,
31'b1000001100000000000000001010000,
31'b1000000010000000000000000000101,
31'b0000100001000000001000100100000,
31'b0000100000010100000000000010000,
31'b0000100000010010000000000010000,
31'b0000100000010000000000000010000,
31'b0001100001000000000000000001000,
31'b0000000000000000000100010000100,
31'b0000100000001010000000000010000,
31'b0000100000001000000000000010000,
31'b0000100000000110000000000010000,
31'b0000100000000100000000000010000,
31'b0000100000000010000000000010000,
31'b0000100000000000000000000010000,
31'b0001100000110000000000000001000,
31'b1100000000000100100000000010000,
31'b0001010000000000100000000000010,
31'b1100000000000000100000000010000,
31'b0010001000000001001000000000100,
31'b1100001000000000001000100000000,
31'b0001010000001000100000000000010,
31'b1100000000001000100000000010000,
31'b0001100000100000000000000001000,
31'b0001000000000101000000000000100,
31'b0000000100000000000000010010000,
31'b0001000000000001000000000000100,
31'b0000100100000000000100000000100,
31'b0001000101000000000000010001000,
31'b0001000001000000010100000000000,
31'b0001000000001001000000000000100,
31'b0001100000010000000000000001000,
31'b0010100011000000000000000100000,
31'b0001100000010100000000000001000,
31'b1100000000100000100000000010000,
31'b0000100000000000001000100100000,
31'b0100000000000101001000000000001,
31'b0100000000000011001000000000001,
31'b0100000000000001001000000000001,
31'b0001100000000000000000000001000,
31'b0001100000000010000000000001000,
31'b0001100000000100000000000001000,
31'b0001000000100001000000000000100,
31'b0000000000000001010000010000000,
31'b0000100001000100000000000010000,
31'b0000100001000010000000000010000,
31'b0000100001000000000000000010000,
31'b1110001100000000000000000000000,
31'b0010100100100000000000000100000,
31'b0001010000000000000100001010000,
31'b1100000000000000000100001000010,
31'b0101000000000000000101000000000,
31'b0110100000010000000000001000000,
31'b0001000000000000101000010000000,
31'b1001000000000000000100000001001,
31'b1010100001000000000010000000000,
31'b0010001000000000100000010000000,
31'b0000010000000000110010000000000,
31'b0010110000000000000001000010000,
31'b0110100000000010000000001000000,
31'b0110100000000000000000001000000,
31'b0001000110000000010100000000000,
31'b1101000100000000001000000000000,
31'b0110000000001000100010000000000,
31'b0010100100000000000000000100000,
31'b1000001010000000000000001010000,
31'b1000000100000000000000000000101,
31'b0110000000000000100010000000000,
31'b0110000000000010100010000000000,
31'b0110000000000100100010000000000,
31'b1000000100001000000000000000101,
31'b0001000010000001000100000010000,
31'b0010100100010000000000000100000,
31'b0000010000000000000000100010001,
31'b1000000100010000000000000000101,
31'b1010001000000000000000001100000,
31'b1010000100000000000010010000000,
31'b1000011100000000010000000000000,
31'b1000000000000000000000101001000,
31'b1000000000000000000100000010001,
31'b1010000000100000100000001000000,
31'b0000000010010000000000010010000,
31'b0100000010000001000000100000010,
31'b0010000000000000000000010100000,
31'b0010000000000010000000010100000,
31'b0000000000000000000110000000010,
31'b0000001000000000000000110001000,
31'b1010100000000000000010000000000,
31'b1010100000000010000010000000000,
31'b0000000010000000000000010010000,
31'b0000001000000001000011000000000,
31'b0010000000010000000000010100000,
31'b0110100001000000000000001000000,
31'b0000000010001000000000010010000,
31'b0000001000010000000000110001000,
31'b1010000000000010100000001000000,
31'b1010000000000000100000001000000,
31'b0100000000010000000010100001000,
31'b1010000000000100100000001000000,
31'b0010000000100000000000010100000,
31'b1010000000001000100000001000000,
31'b0100000000000001000001010000000,
31'b0100001010000000000010000010000,
31'b1010100000100000000010000000000,
31'b1010000000010000100000001000000,
31'b0100000000000000000010100001000,
31'b0100001000000000000100010000010,
31'b0010101100000000100000000000000,
31'b0001010000000000000000100001001,
31'b0100000000010001000001010000000,
31'b0000000010000001000100000001000,
31'b0000100001000000000000000100011,
31'b0000100000010001010000000000000,
31'b0000000001010000000000010010000,
31'b0100100000000000000000001110000,
31'b0110010000000000000000000001100,
31'b0001000000010000000000010001000,
31'b0001000100010000010100000000000,
31'b0001000100000000100001000000001,
31'b0000100000000011010000000000000,
31'b0000100000000001010000000000000,
31'b0000000001000000000000010010000,
31'b0000100000000101010000000000000,
31'b0001000000000010000000010001000,
31'b0001000000000000000000010001000,
31'b0001000100000000010100000000000,
31'b0001000000000100000000010001000,
31'b1100000000000000100100000000100,
31'b0010100110000000000000000100000,
31'b1000001000000000000000001010000,
31'b1000001000000010000000001010000,
31'b1100011000000000000001000000000,
31'b0001001000000000000001000010010,
31'b1000110000000000000000100000100,
31'b0000100100010000000000000010000,
31'b0001000000000001000100000010000,
31'b0000100000100001010000000000000,
31'b0000000000000000010000000001100,
31'b0000100100001000000000000010000,
31'b0001000000100010000000010001000,
31'b0001000000100000000000010001000,
31'b0000100100000010000000000010000,
31'b0000100100000000000000000010000,
31'b0000100000000000000000000100011,
31'b0100000000000101000000100000010,
31'b0000000000010000000000010010000,
31'b0100000000000001000000100000010,
31'b0010000010000000000000010100000,
31'b0011000000000000000001001000100,
31'b0000000010000000000110000000010,
31'b0100001000100000000010000010000,
31'b0000000000000100000000010010000,
31'b0000100001000001010000000000000,
31'b0000000000000000000000010010000,
31'b0000000000000010000000010010000,
31'b0000100000000000000100000000100,
31'b0001000001000000000000010001000,
31'b0000000000001000000000010010000,
31'b0000000000100001000100000001000,
31'b0001100100010000000000000001000,
31'b1100001000000000000000000000011,
31'b0000001000000000000001000001010,
31'b0100001000001000000010000010000,
31'b0010000010100000000000010100000,
31'b1100000000000001110000000000000,
31'b0100001000000010000010000010000,
31'b0100001000000000000010000010000,
31'b0001100100000000000000000001000,
31'b0001100100000010000000000001000,
31'b0000000000100000000000010010000,
31'b0000000000100010000000010010000,
31'b0000100000100000000100000000100,
31'b0001000000000000010000000010100,
31'b0000000000101000000000010010000,
31'b0000000000000001000100000001000,
31'b1110010000000000000000000000000,
31'b0011000000000000000000000010010,
31'b1110010000000100000000000000000,
31'b0011000000000100000000000010010,
31'b1110010000001000000000000000000,
31'b0011000000001000000000000010010,
31'b1000000000110000010000000000000,
31'b1011000000000000000010000000001,
31'b0000000000000000100000100000010,
31'b1001000000000000000000010000100,
31'b1000000000101000010000000000000,
31'b1001000000000100000000010000100,
31'b1000000000100100010000000000000,
31'b1001000000001000000000010000100,
31'b1000000000100000010000000000000,
31'b1000000000100010010000000000000,
31'b1110010000100000000000000000000,
31'b0011000000100000000000000010010,
31'b1000000000011000010000000000000,
31'b1000011000000000000000000000101,
31'b1000000000010100010000000000000,
31'b1100000000000000001000010000001,
31'b1000000000010000010000000000000,
31'b1000000000010010010000000000000,
31'b1000000000001100010000000000000,
31'b1001000000100000000000010000100,
31'b1000000000001000010000000000000,
31'b1000000000001010010000000000000,
31'b1000000000000100010000000000000,
31'b1000000000000110010000000000000,
31'b1000000000000000010000000000000,
31'b1000000000000010010000000000000,
31'b1110010001000000000000000000000,
31'b0011000001000000000000000010010,
31'b0100100000000000110000000000000,
31'b0110000000000000000011000010000,
31'b0010000000000100000000000001010,
31'b0010010000000000000010001000000,
31'b0010000000000000000000000001010,
31'b0010000000000010000000000001010,
31'b1000100000000000000100000001000,
31'b1001000001000000000000010000100,
31'b1000100000000100000100000001000,
31'b1000100100000000010000010000000,
31'b1000100000001000000100000001000,
31'b0100001000000000001000001000001,
31'b1000000001100000010000000000000,
31'b1001000100000001000000000001000,
31'b0001001000000010000000001000100,
31'b0001001000000000000000001000100,
31'b1000010000000000100100000000010,
31'b1000001000000000110000000100000,
31'b1100100000000000000000100000010,
31'b0010100000000001000000000000110,
31'b1000000001010000010000000000000,
31'b1000000001010010010000000000000,
31'b1000100000100000000100000001000,
31'b1001000000000000010000000011000,
31'b1000000001001000010000000000000,
31'b1000000000000001000100000000100,
31'b1000000001000100010000000000000,
31'b1000100000000001000000010010000,
31'b1000000001000000010000000000000,
31'b1000000001000010010000000000000,
31'b1110010010000000000000000000000,
31'b0011000010000000000000000010010,
31'b0001001001000000100000000000010,
31'b0001000000000000000100000000101,
31'b1100000100100000000001000000000,
31'b0001100000000000000000010010001,
31'b1010000100000001000000000100000,
31'b0001000000010000000000000100010,
31'b1000000000000000000001001100000,
31'b1001000010000000000000010000100,
31'b1000000010101000010000000000000,
31'b0001000000001000000000000100010,
31'b1000000010100100010000000000000,
31'b0001000000000100000000000100010,
31'b1000000010100000010000000000000,
31'b0001000000000000000000000100010,
31'b1100000100001000000001000000000,
31'b0000000101000000000011001000000,
31'b1000010100000000000000001010000,
31'b0000000100001000000000000001001,
31'b1100000100000000000001000000000,
31'b0000000100000100000000000001001,
31'b1000000010010000010000000000000,
31'b0000000100000000000000000001001,
31'b1000000010001100010000000000000,
31'b0000000000001000100001010000000,
31'b1000000010001000010000000000000,
31'b0000000000000000000000101000100,
31'b1000000010000100010000000000000,
31'b0000000000000000100001010000000,
31'b1000000010000000010000000000000,
31'b0100000000000000001100000000000,
31'b0001001000000100100000000000010,
31'b1100100000000000000001010000000,
31'b0001001000000000100000000000010,
31'b1000100000000000101100000000000,
31'b0010010000000001001000000000100,
31'b1100010000000000001000100000000,
31'b0010000010000000000000000001010,
31'b0010000010000010000000000001010,
31'b0000100100000000100001000000000,
31'b0100100000000000011000000001000,
31'b0001010000000000000001000100001,
31'b0010001000000000000000100010010,
31'b0100000100000000001000000010100,
31'b0100000000000000000011000100000,
31'b1000000011100000010000000000000,
31'b0010000000100001000010000000000,
31'b0001000100000000000000000010001,
31'b0000000100000000000011001000000,
31'b0001001000100000100000000000010,
31'b0010000000011001000010000000000,
31'b1100000101000000000001000000000,
31'b0010000000010101000010000000000,
31'b1001000100000000000010000000010,
31'b0010000000010001000010000000000,
31'b0001111000000000000000000001000,
31'b0010000100000000100000100000001,
31'b1000000011001000010000000000000,
31'b0010000000001001000010000000000,
31'b1000101000000000000011000000000,
31'b0010000000000101000010000000000,
31'b1000000011000000010000000000000,
31'b0010000000000001000010000000000,
31'b1000000000010001000000000010000,
31'b1100000000000000000000110000010,
31'b1100000000000000010000001100000,
31'b0000101000100000010000001000000,
31'b1100000010100000000001000000000,
31'b0000101010000000000001000100000,
31'b1010000010000001000000000100000,
31'b0000000010100000000000000001001,
31'b1000000000000001000000000010000,
31'b1000000000000011000000000010000,
31'b1000000000000101000000000010000,
31'b1000100001000000010000010000000,
31'b1000000000001001000000000010000,
31'b1000000000100000000100010001000,
31'b1000000100100000010000000000000,
31'b1001000001000001000000000001000,
31'b1100000010001000000001000000000,
31'b0000101000000100010000001000000,
31'b1000010010000000000000001010000,
31'b0000101000000000010000001000000,
31'b1100000010000000000001000000000,
31'b0000000010000100000000000001001,
31'b1000000100010000010000000000000,
31'b0000000010000000000000000001001,
31'b1000000000100001000000000010000,
31'b1000000000100011000000000010000,
31'b1000000100001000010000000000000,
31'b1000100000000000000000000011100,
31'b0000000000000000101000000000001,
31'b1000000000000000000100010001000,
31'b1000000100000000010000000000000,
31'b1000000100000010010000000000000,
31'b1100100000000000001000000000001,
31'b0000100010000000010100000000001,
31'b0110000000000000001000000100100,
31'b0000100000000000001001000001000,
31'b0010011000000000000000010100000,
31'b0000001000000000000100001001000,
31'b0010000100000000000000000001010,
31'b0000000000000000010010000100000,
31'b1000000001000001000000000010000,
31'b1000100000000100010000010000000,
31'b1000100000000010010000010000000,
31'b1000100000000000010000010000000,
31'b1001100000100000000000000000100,
31'b1001000000000101000000000001000,
31'b1001000000000011000000000001000,
31'b1001000000000001000000000001000,
31'b0001000010000000000000000010001,
31'b0000001000000000001000000100001,
31'b0011000000000000000100000000110,
31'b0000101001000000010000001000000,
31'b1100000011000000000001000000000,
31'b0000001000100000000100001001000,
31'b1001000010000000000010000000010,
31'b0000000011000000000000000001001,
31'b1001100000001000000000000000100,
31'b0110010000000000000010000100000,
31'b1001000000000000000100010010000,
31'b1000100000100000010000010000000,
31'b1001100000000000000000000000100,
31'b1001100000000010000000000000100,
31'b1000000101000000010000000000000,
31'b1001000000100001000000000001000,
31'b1100000000101000000001000000000,
31'b0000101000001000000001000100000,
31'b1010000000001001000000000100000,
31'b0000000000101000000000000001001,
31'b1100000000100000000001000000000,
31'b0000101000000000000001000100000,
31'b1010000000000001000000000100000,
31'b0000000000100000000000000001001,
31'b1000000010000001000000000010000,
31'b1000001000000000000011010000000,
31'b1010010000000000010001000000000,
31'b0101000000000000001000000001100,
31'b1100000000110000000001000000000,
31'b0001011000000000000000010001000,
31'b1010000000010001000000000100000,
31'b0001000100000000000000000100010,
31'b1100000000001000000001000000000,
31'b0000000001000000000011001000000,
31'b1000010000000000000000001010000,
31'b0000000000001000000000000001001,
31'b1100000000000000000001000000000,
31'b0000000000000100000000000001001,
31'b0000000000000010000000000001001,
31'b0000000000000000000000000001001,
31'b1100000000011000000001000000000,
31'b0010000001000000100000100000001,
31'b1000010000010000000000001010000,
31'b0000000100000000000000101000100,
31'b1100000000010000000001000000000,
31'b0000000100000000100001010000000,
31'b1000000110000000010000000000000,
31'b0000000000010000000000000001001,
31'b0001000000100000000000000010001,
31'b0000100000000000010100000000001,
31'b0001001100000000100000000000010,
31'b0000100010000000001001000001000,
31'b1100000001100000000001000000000,
31'b0000101001000000000001000100000,
31'b1010000001000001000000000100000,
31'b0000000010000000010010000100000,
31'b0000100000000000100001000000000,
31'b0010000000000000010010000010000,
31'b0000100000000100100001000000000,
31'b1010001000000001100000000000000,
31'b0100000000000000001000000010100,
31'b0100000100000000000011000100000,
31'b0100010000000000000101100000000,
31'b1010000000000000010000000000011,
31'b0001000000000000000000000010001,
31'b0000000000000000000011001000000,
31'b0001000000000100000000000010001,
31'b0000000001001000000000000001001,
31'b1100000001000000000001000000000,
31'b0000000001000100000000000001001,
31'b1001000000000000000010000000010,
31'b0000000001000000000000000001001,
31'b0001000000010000000000000010001,
31'b0010000000000000100000100000001,
31'b0001100000000000000000010100010,
31'b0010000100001001000010000000000,
31'b1100000001010000000001000000000,
31'b0010000100000101000010000000000,
31'b1001000000010000000010000000010,
31'b0010000100000001000010000000000,
31'b1110011000000000000000000000000,
31'b0011001000000000000000000010010,
31'b0001000100000000000100001010000,
31'b1100000000000000010010010000000,
31'b0000100000000011000000001010000,
31'b0000100000000001000000001010000,
31'b0000000001000000010000011000000,
31'b0100100000010000010000000100000,
31'b1000000000000000001010000000001,
31'b1001001000000000000000010000100,
31'b0000000100000000110010000000000,
31'b0100100000001000010000000100000,
31'b0000000000000100001000000010010,
31'b0100100000000100010000000100000,
31'b0000000000000000001000000010010,
31'b0100100000000000010000000100000,
31'b0111000010000000000100000000000,
31'b0010110000000000000000000100000,
31'b1000010000000010000000000000101,
31'b1000010000000000000000000000101,
31'b1101000000000000000010000000100,
31'b0011000000000001000010100000000,
31'b1000001000010000010000000000000,
31'b1000010000001000000000000000101,
31'b1000001000001100010000000000000,
31'b0100100010000000000001001000000,
31'b1000001000001000010000000000000,
31'b1000010000010000000000000000101,
31'b1000001000000100010000000000000,
31'b1010010000000000000010010000000,
31'b1000001000000000010000000000000,
31'b1000001000000010010000000000000,
31'b0001000010000100100000000000010,
31'b0001000000100000000000001000100,
31'b0001000010000000100000000000010,
31'b1000000010000000000000110000100,
31'b0000000000000100010000011000000,
31'b0000000000000000000000100100010,
31'b0000000000000000010000011000000,
31'b0000000000000100000000100100010,
31'b1000101000000000000100000001000,
31'b0001000000000000001000000001010,
31'b0001010000000000001010001000000,
31'b0010000010000000000000100010010,
31'b0100000000000010001000001000001,
31'b0100000000000000001000001000001,
31'b0000000001000000001000000010010,
31'b0100100001000000010000000100000,
31'b0001000000000010000000001000100,
31'b0001000000000000000000001000100,
31'b1000000000001000000001000000110,
31'b1000000000000000110000000100000,
31'b1001000010000000010000100000000,
31'b0001000000001000000000001000100,
31'b1000000000000000000001000000110,
31'b1000000000001000110000000100000,
31'b0110010000000000000000011000000,
31'b0100000000000000000100000101000,
31'b1000001001001000010000000000000,
31'b1000001000000001000100000000100,
31'b1000100010000000000011000000000,
31'b0100000000100000001000001000001,
31'b1000001001000000010000000000000,
31'b1000010000000001100001000000000,
31'b0100000000000000100011000000000,
31'b0110100000000000010000000010000,
31'b0001000001000000100000000000010,
31'b1000000001000000000000110000100,
31'b0110000100000000000000000001100,
31'b0000100100000000000001000100000,
31'b0001010000010000010100000000000,
31'b0001010000000000100001000000001,
31'b1000001000000000000001001100000,
31'b1000000100000000000011010000000,
31'b0001010000001000010100000000000,
31'b0010100000000001000000001100000,
31'b0011000000000000000000100001010,
31'b0001010100000000000000010001000,
31'b0001010000000000010100000000000,
31'b0001001000000000000000000100010,
31'b0111000000000000000100000000000,
31'b0111000000000010000100000000000,
31'b0111000000000100000100000000000,
31'b1000010010000000000000000000101,
31'b1100001100000000000001000000000,
31'b0000110000010100000000000010000,
31'b1000100100000000000000100000100,
31'b0000110000010000000000000010000,
31'b0111000000010000000100000000000,
31'b0100100000000000000001001000000,
31'b1000100000000000000000001001001,
31'b0000110000001000000000000010000,
31'b1000100001000000000011000000000,
31'b0000110000000100000000000010000,
31'b1000001010000000010000000000000,
31'b0000110000000000000000000010000,
31'b0001000000000100100000000000010,
31'b1000000000001000100001001000000,
31'b0001000000000000100000000000010,
31'b1000000000000000000000110000100,
31'b1001000000100000010000100000000,
31'b1000000000000000100001001000000,
31'b0001000000001000100000000000010,
31'b1000000000001000000000110000100,
31'b0001110000100000000000000001000,
31'b0010000000000100000000100010010,
31'b0001000000010000100000000000010,
31'b0010000000000000000000100010010,
31'b1000100000100000000011000000000,
31'b1010000000000000000010100000001,
31'b0001010001000000010100000000000,
31'b0010001000100001000010000000000,
31'b0000000000000000000001010100000,
31'b0001000010000000000000001000100,
31'b0001000000100000100000000000010,
31'b1000000010000000110000000100000,
31'b1001000000000000010000100000000,
31'b1001000000000010010000100000000,
31'b1001000000000100010000100000000,
31'b0110000000000000000100000011000,
31'b0001110000000000000000000001000,
31'b0100100001000000000001001000000,
31'b0001110000000100000000000001000,
31'b0010001000001001000010000000000,
31'b1000100000000000000011000000000,
31'b1010000000000000110000000010000,
31'b1000100000000100000011000000000,
31'b0010001000000001000010000000000,
31'b1100000000000000000110000001000,
31'b0000100010001000000001000100000,
31'b0001000000000000000100001010000,
31'b0000100000100000010000001000000,
31'b0110000010000000000000000001100,
31'b0000100010000000000001000100000,
31'b0001010000000000101000010000000,
31'b0000100010000100000001000100000,
31'b1000001000000001000000000010000,
31'b1000001000000011000000000010000,
31'b0000000000000000110010000000000,
31'b0010100000000000000001000010000,
31'b1000001000001001000000000010000,
31'b0110110000000000000000001000000,
31'b0000000100000000001000000010010,
31'b0110000000000000101000000000100,
31'b0000100000000110010000001000000,
31'b0000100000000100010000001000000,
31'b0000100000000010010000001000000,
31'b0000100000000000010000001000000,
31'b1100001010000000000001000000000,
31'b0000100010100000000001000100000,
31'b1000100010000000000000100000100,
31'b0000100000001000010000001000000,
31'b0000000000000100000000100010001,
31'b0100100000000001000000000110000,
31'b0000000000000000000000100010001,
31'b0000100000010000010000001000000,
31'b1000000000000000000010100000010,
31'b1000001000000000000100010001000,
31'b1000001100000000010000000000000,
31'b1000010000000000000000101001000,
31'b1010000000000001001000000001000,
31'b0000000000100000001000000100001,
31'b0001000110000000100000000000010,
31'b0000101000000000001001000001000,
31'b0010010000000000000000010100000,
31'b0000000000000000000100001001000,
31'b0000010000000000000110000000010,
31'b0000001000000000010010000100000,
31'b1010110000000000000010000000000,
31'b0101000000001000000000000100100,
31'b0000010010000000000000010010000,
31'b1010000010000001100000000000000,
31'b0101000000000010000000000100100,
31'b0101000000000000000000000100100,
31'b0000010010001000000000010010000,
31'b1100000000000000110000001000000,
31'b0000000000000010001000000100001,
31'b0000000000000000001000000100001,
31'b0100100000000001001000100000000,
31'b0000100001000000010000001000000,
31'b0010010000100000000000010100000,
31'b0000000000100000000100001001000,
31'b1100100000000000010010000000000,
31'b0000100010000000001110000000000,
31'b0100000000000100010000010100000,
31'b0100000000000000000000101000010,
31'b0100000000000000010000010100000,
31'b0100000000000100000000101000010,
31'b1001101000000000000000000000100,
31'b0001000000000000000000100001001,
31'b1101000000000000000001100000000,
31'b0011000000000001000001000000100,
31'b0110000000001000000000000001100,
31'b0000100000001000000001000100000,
31'b0001000101000000100000000000010,
31'b0000100010100000010000001000000,
31'b0110000000000000000000000001100,
31'b0000100000000000000001000100000,
31'b1010001000000001000000000100000,
31'b0000100000000100000001000100000,
31'b1000001010000001000000000010000,
31'b1000000000000000000011010000000,
31'b0000010001000000000000010010000,
31'b1010000001000001100000000000000,
31'b0110000000010000000000000001100,
31'b0001010000000000000000010001000,
31'b0001010100000000010100000000000,
31'b0001010000000100000000010001000,
31'b1100001000001000000001000000000,
31'b0000100010000100010000001000000,
31'b1000100000001000000000100000100,
31'b0000100010000000010000001000000,
31'b1100001000000000000001000000000,
31'b0000100000100000000001000100000,
31'b1000100000000000000000100000100,
31'b0000001000000000000000000001001,
31'b0011000000000000001000000001001,
31'b1100000000000001000100000000010,
31'b0000010000000000010000000001100,
31'b0000110100001000000000000010000,
31'b1100001000010000000001000000000,
31'b0001010000100000000000010001000,
31'b1000100000010000000000100000100,
31'b0000110100000000000000000010000,
31'b0001001000100000000000000010001,
31'b0000101000000000010100000000001,
31'b0001000100000000100000000000010,
31'b1010000000010001100000000000000,
31'b0110000001000000000000000001100,
31'b0000100001000000000001000100000,
31'b0001000100001000100000000000010,
31'b0000100001000100000001000100000,
31'b0000101000000000100001000000000,
31'b1010000000000101100000000000000,
31'b0000010000000000000000010010000,
31'b1010000000000001100000000000000,
31'b0100000000000000000001011000000,
31'b0101000010000000000000000100100,
31'b0000010000001000000000010010000,
31'b1010000000001001100000000000000,
31'b0001001000000000000000000010001,
31'b0000001000000000000011001000000,
31'b0001001000000100000000000010001,
31'b0000100011000000010000001000000,
31'b1100001001000000000001000000000,
31'b0000100001100000000001000100000,
31'b1001001000000000000010000000010,
31'b0000100000000000001110000000000,
31'b0001110100000000000000000001000,
31'b1100000000000000100001000100000,
31'b0000010000100000000000010010000,
31'b1010000000100001100000000000000,
31'b1100000000000000010000000000110,
31'b0010000000000100001000000010001,
31'b0010000000000010001000000010001,
31'b0010000000000000001000000010001,
31'b1110100000000000000000000000000,
31'b0010001000100000000000000100000,
31'b0000000000100000000000100001000,
31'b0100001000000001000001000000000,
31'b1110100000001000000000000000000,
31'b0010100001000000000010001000000,
31'b0100000000010000000100000000010,
31'b0100001000001001000001000000000,
31'b1110100000010000000000000000000,
31'b0010100100000000100000010000000,
31'b0100000000001000000100000000010,
31'b0100001000010001000001000000000,
31'b0100000000000100000100000000010,
31'b0110001100000000000000001000000,
31'b0100000000000000000100000000010,
31'b0100000000000010000100000000010,
31'b0000000000000100000000100001000,
31'b0010001000000000000000000100000,
31'b0000000000000000000000100001000,
31'b0000000000000010000000100001000,
31'b0010000001010000100000000000000,
31'b0010001000001000000000000100000,
31'b0000000000001000000000100001000,
31'b0000001010010000000000000010000,
31'b0010000001001000100000000000000,
31'b0010001000010000000000000100000,
31'b0000000000010000000000100001000,
31'b0000001010001000000000000010000,
31'b0010000001000000100000000000000,
31'b0010000001000010100000000000000,
31'b0001000000000000001000000100000,
31'b0000001010000000000000000010000,
31'b1110100001000000000000000000000,
31'b0010100000001000000010001000000,
31'b0100010000000000110000000000000,
31'b0100010000000010110000000000000,
31'b0010000000110000100000000000000,
31'b0010100000000000000010001000000,
31'b0100010000001000110000000000000,
31'b1001000100000000001010000000000,
31'b1000010000000000000100000001000,
31'b1010000000000000000000011100000,
31'b1010000000000000010000100000010,
31'b1000010100000000010000010000000,
31'b0010000000100000100000000000000,
31'b0010000000100010100000000000000,
31'b0100000001000000000100000000010,
31'b0100001000000000100000000000101,
31'b0010000000011000100000000000000,
31'b0010001001000000000000000100000,
31'b0000000001000000000000100001000,
31'b0001001000000000101000000000000,
31'b0010000000010000100000000000000,
31'b0001000000000000000000100010000,
31'b0010000000010100100000000000000,
31'b0010000010000000001000000001000,
31'b0010000000001000100000000000000,
31'b0010000000001010100000000000000,
31'b0010000000001100100000000000000,
31'b0011000010000000000000100100000,
31'b0010000000000000100000000000000,
31'b0010000000000010100000000000000,
31'b0010000000000100100000000000000,
31'b0010000000000110100000000000000,
31'b1110100010000000000000000000000,
31'b0010100000000000011100000000000,
31'b0100000000000000000010010010000,
31'b0100001010000001000001000000000,
31'b1100000000000000000000010000011,
31'b0001010000000000000000010010001,
31'b0100000010010000000100000000010,
31'b0000001000110000000000000010000,
31'b0001001001100000000000000001000,
31'b0000001100000001010000000000000,
31'b0100000010001000000100000000010,
31'b0000001000101000000000000010000,
31'b0110000000000000000000000010101,
31'b0000001000100100000000000010000,
31'b0100000010000000000100000000010,
31'b0000001000100000000000000010000,
31'b0011000000000000001000000010000,
31'b0010001010000000000000000100000,
31'b0000000010000000000000100001000,
31'b0000001000011000000000000010000,
31'b0011000000001000001000000010000,
31'b0001000000000000100000000101000,
31'b0000001000010010000000000010000,
31'b0000001000010000000000000010000,
31'b0001001001000000000000000001000,
31'b0000000000000000101000100000000,
31'b0000001000001010000000000010000,
31'b0000001000001000000000000010000,
31'b0010000011000000100000000000000,
31'b0000001000000100000000000010000,
31'b0000001000000010000000000010000,
31'b0000001000000000000000000010000,
31'b0001001000110000000000000001000,
31'b1100010000000000000001010000000,
31'b0000010000000000000000010001001,
31'b1000010000000000101100000000000,
31'b0010100000000001001000000000100,
31'b1100100000000000001000100000000,
31'b1000000000000010000000011010000,
31'b1000000000000000000000011010000,
31'b0001001000100000000000000001000,
31'b0101000000000001000001100000000,
31'b0001100000000000000001000100001,
31'b0011000000100000000000100100000,
31'b0010000010100000100000000000000,
31'b0010000010100010100000000000000,
31'b0100000100000000100000001010000,
31'b0010000000000000000000001000110,
31'b0001001000010000000000000001000,
31'b0010001011000000000000000100000,
31'b0000000000000000100000000110000,
31'b0010000000001000001000000001000,
31'b0010000010010000100000000000000,
31'b0010000000000100001000000001000,
31'b0010000000000010001000000001000,
31'b0010000000000000001000000001000,
31'b0001001000000000000000000001000,
31'b0001001000000010000000000001000,
31'b0001001000000100000000000001000,
31'b0011000000000000000000100100000,
31'b0010000010000000100000000000000,
31'b0010000010000010100000000000000,
31'b0010000010000100100000000000000,
31'b0000001001000000000000000010000,
31'b1110100100000000000000000000000,
31'b0010100000010000100000010000000,
31'b0101000000000000001000001000000,
31'b0101000000000010001000001000000,
31'b0001010000000000001001000010000,
31'b1100000000000000001001000000010,
31'b0001000000000000000100100000100,
31'b1001000001000000001010000000000,
31'b1010001001000000000010000000000,
31'b0010100000000000100000010000000,
31'b0101000000010000001000001000000,
31'b1000010001000000010000010000000,
31'b0110001000000010000000001000000,
31'b0110001000000000000000001000000,
31'b0100000100000000000100000000010,
31'b0110001000000100000000001000000,
31'b0010000000000000000010011000000,
31'b0010001100000000000000000100000,
31'b0000000100000000000000100001000,
31'b0000011000000000010000001000000,
31'b0010000101010000100000000000000,
31'b1110000001000000000000010000000,
31'b0000000100001000000000100001000,
31'b0000110010000000000000000001001,
31'b0010000101001000100000000000000,
31'b0010100000100000100000010000000,
31'b0000000100010000000000100001000,
31'b1000010000000000000000000011100,
31'b0010000101000000100000000000000,
31'b0110001000100000000000001000000,
31'b0000000000000000000000001000101,
31'b0000001110000000000000000010000,
31'b1100010000000000001000000000001,
31'b0001000000000101010000100000000,
31'b0101000001000000001000001000000,
31'b0001000000000001010000100000000,
31'b0010101000000000000000010100000,
31'b1110000000100000000000010000000,
31'b1001000000000010001010000000000,
31'b1001000000000000001010000000000,
31'b1010001000000000000010000000000,
31'b1010001000000010000010000000000,
31'b1010001000000100000010000000000,
31'b1000010000000000010000010000000,
31'b0010000100100000100000000000000,
31'b0110001001000000000000001000000,
31'b0100000101000000000100000000010,
31'b1001000000010000001010000000000,
31'b0010000100011000100000000000000,
31'b1110000000001000000000010000000,
31'b0000000101000000000000100001000,
31'b0001001100000000101000000000000,
31'b0010000100010000100000000000000,
31'b1110000000000000000000010000000,
31'b0010000100010100100000000000000,
31'b1110000000000100000000010000000,
31'b0010000100001000100000000000000,
31'b0110100000000000000010000100000,
31'b0010000100001100100000000000000,
31'b1100000000000000000010000000101,
31'b0010000100000000100000000000000,
31'b0100000000000000000000000010110,
31'b0010000100000100100000000000000,
31'b0110000010000000000100000000001,
31'b0000010001010000100001000000000,
31'b0000001000010001010000000000000,
31'b1011000000000000000010100000000,
31'b1001000000000000010100001000000,
31'b0000010000000001000000000000101,
31'b0000011000000000000001000100000,
31'b0011000000000001011000000000000,
31'b0000110000100000000000000001001,
31'b0000010001000000100001000000000,
31'b0000001000000001010000000000000,
31'b1010100000000000010001000000000,
31'b1000000000000000100010000010000,
31'b0000001001000000000100000000100,
31'b0000000000000000100000000000011,
31'b0100000110000000000100000000010,
31'b0000001100100000000000000010000,
31'b1100000000000000001000110000000,
31'b0010001110000000000000000100000,
31'b1000100000000000000000001010000,
31'b1000100000000010000000001010000,
31'b1100110000000000000001000000000,
31'b0001100000000000000001000010010,
31'b1000100000001000000000001010000,
31'b0000110000000000000000000001001,
31'b0101010000000001001000000000000,
31'b0000001000100001010000000000000,
31'b1000100000010000000000001010000,
31'b1000000000000000010000100000001,
31'b0010000111000000100000000000000,
31'b0000001100000100000000000010000,
31'b0000001100000010000000000010000,
31'b0000001100000000000000000010000,
31'b0000010000010000100001000000000,
31'b0000010000000000010100000000001,
31'b0000101000010000000000010010000,
31'b0011000000000000001100000000100,
31'b0000001000010000000100000000100,
31'b0000011001000000000001000100000,
31'b1001000000000001000000001000100,
31'b1001000010000000001010000000000,
31'b0000010000000000100001000000000,
31'b0000010000000010100001000000000,
31'b0000101000000000000000010010000,
31'b1000010010000000010000010000000,
31'b0000001000000000000100000000100,
31'b0000001000000010000100000000100,
31'b0100000000000000100000001010000,
31'b0110000000100000000100000000001,
31'b0001110000000000000000000010001,
31'b1100100000000000000000000000011,
31'b0000100000000000000001000001010,
31'b0110000000000000000000000100110,
31'b0010000110010000100000000000000,
31'b1110000010000000000000010000000,
31'b0110000000000000110001000000000,
31'b0100100000000000000010000010000,
31'b0001001100000000000000000001000,
31'b0001010000000000010000101000000,
31'b0001010000000000000000010100010,
31'b1100000000000000000000010110000,
31'b0010000110000000100000000000000,
31'b0110000000000100000100000000001,
31'b0110000000000010000100000000001,
31'b0110000000000000000100000000001,
31'b1000000000000001000000000001001,
31'b0010000000100000000000000100000,
31'b0100000000000011000001000000000,
31'b0100000000000001000001000000000,
31'b1010000000000000100000011000000,
31'b0010000000101000000000000100000,
31'b0100001000010000000100000000010,
31'b0100000000001001000001000000000,
31'b1010000101000000000010000000000,
31'b0010000000110000000000000100000,
31'b0100001000001000000100000000010,
31'b0100000000010001000001000000000,
31'b0110000100000010000000001000000,
31'b0110000100000000000000001000000,
31'b0100001000000000000100000000010,
31'b0000000010100000000000000010000,
31'b0010000000000010000000000100000,
31'b0010000000000000000000000100000,
31'b0000001000000000000000100001000,
31'b0010000000000100000000000100000,
31'b0010000000001010000000000100000,
31'b0010000000001000000000000100000,
31'b0000001000001000000000100001000,
31'b0000000010010000000000000010000,
31'b0010000000010010000000000100000,
31'b0010000000010000000000000100000,
31'b0000001000010000000000100001000,
31'b0000000010001000000000000010000,
31'b0010001001000000100000000000000,
31'b0000000010000100000000000010000,
31'b0000000010000010000000000010000,
31'b0000000010000000000000000010000,
31'b1010000100010000000010000000000,
31'b0010000001100000000000000100000,
31'b0100011000000000110000000000000,
31'b0100000001000001000001000000000,
31'b0010100100000000000000010100000,
31'b0010101000000000000010001000000,
31'b1000000100000000000000010000101,
31'b1001000000000001000000000010001,
31'b1010000100000000000010000000000,
31'b1010000100000010000010000000000,
31'b1010000100000100000010000000000,
31'b0100000001010001000001000000000,
31'b0010001000100000100000000000000,
31'b0110000101000000000000001000000,
31'b0100001001000000000100000000010,
31'b0100000000000000100000000000101,
31'b0010000001000010000000000100000,
31'b0010000001000000000000000100000,
31'b0001000000000010101000000000000,
31'b0001000000000000101000000000000,
31'b0010001000010000100000000000000,
31'b0010000001001000000000000100000,
31'b0011000000000000000000000111000,
31'b0001000000001000101000000000000,
31'b0001000010000000000000000001000,
31'b0010000001010000000000000100000,
31'b0010000000000000001000100010000,
31'b0001000000010000101000000000000,
31'b0010001000000000100000000000000,
31'b0010001000000010100000000000000,
31'b0010001000000100100000000000000,
31'b0000000011000000000000000010000,
31'b1011000000000000010000000000010,
31'b0010000010100000000000000100000,
31'b0100001000000000000010010010000,
31'b0100000010000001000001000000000,
31'b0000010100000010000001000100000,
31'b0000010100000000000001000100000,
31'b0000000000110010000000000010000,
31'b0000000000110000000000000010000,
31'b0001000001100000000000000001000,
31'b0000000100000001010000000000000,
31'b0000000000101010000000000010000,
31'b0000000000101000000000000010000,
31'b0000000101000000000100000000100,
31'b0000000000100100000000000010000,
31'b0000000000100010000000000010000,
31'b0000000000100000000000000010000,
31'b0010000010000010000000000100000,
31'b0010000010000000000000000100000,
31'b0000001010000000000000100001000,
31'b0000000000011000000000000010000,
31'b0000000001000000001000100100000,
31'b0000000000010100000000000010000,
31'b0000000000010010000000000010000,
31'b0000000000010000000000000010000,
31'b0001000001000000000000000001000,
31'b0000000000001100000000000010000,
31'b0000000000001010000000000010000,
31'b0000000000001000000000000010000,
31'b0000000000000110000000000010000,
31'b0000000000000100000000000010000,
31'b0000000000000010000000000010000,
31'b0000000000000000000000000010000,
31'b0001000000110000000000000001000,
31'b0010000011100000000000000100000,
31'b0001110000000000100000000000010,
31'b1100100000000000100000000010000,
31'b0000000100010000000100000000100,
31'b1000010000000000000100100010000,
31'b1000000100000000000010000110000,
31'b1000000000000000001001000000100,
31'b0001000000100000000000000001000,
31'b0001000000100010000000000001000,
31'b0001000000100100000000000001000,
31'b0001100000000001000000000000100,
31'b0000000100000000000100000000100,
31'b0000000100000010000100000000100,
31'b0000000100000100000100000000100,
31'b0000000001100000000000000010000,
31'b0001000000010000000000000001000,
31'b0010000011000000000000000100000,
31'b0001000000010100000000000001000,
31'b0001000010000000101000000000000,
31'b0000000000000000001000100100000,
31'b0000000001010100000000000010000,
31'b0000000001010010000000000010000,
31'b0000000001010000000000000010000,
31'b0001000000000000000000000001000,
31'b0001000000000010000000000001000,
31'b0001000000000100000000000001000,
31'b0000000001001000000000000010000,
31'b0001000000001000000000000001000,
31'b0000000001000100000000000010000,
31'b0000000001000010000000000010000,
31'b0000000001000000000000000010000,
31'b1010000001010000000010000000000,
31'b0010000100100000000000000100000,
31'b0101001000000000001000001000000,
31'b0100000100000001000001000000000,
31'b0110000000010010000000001000000,
31'b0110000000010000000000001000000,
31'b1000000001000000000000010000101,
31'b0110000000010100000000001000000,
31'b1010000001000000000010000000000,
31'b0000000010000001010000000000000,
31'b1010000001000100000010000000000,
31'b0010010000000000000001000010000,
31'b0110000000000010000000001000000,
31'b0110000000000000000000001000000,
31'b0110000000000110000000001000000,
31'b0110000000000100000000001000000,
31'b0010000100000010000000000100000,
31'b0010000100000000000000000100000,
31'b0000010000000010010000001000000,
31'b0000010000000000010000001000000,
31'b0110100000000000100010000000000,
31'b0100000000000000010001000010000,
31'b1000010010000000000000100000100,
31'b0000010000001000010000001000000,
31'b1010000001100000000010000000000,
31'b0010000100010000000000000100000,
31'b0000110000000000000000100010001,
31'b0000010000010000010000001000000,
31'b0110000000100010000000001000000,
31'b0110000000100000000000001000000,
31'b0000001000000000000000001000101,
31'b0000000110000000000000000010000,
31'b1010000000010000000010000000000,
31'b1010000000010010000010000000000,
31'b1010000000010100000010000000000,
31'b0100000101000001000001000000000,
31'b0010100000000000000000010100000,
31'b0110000001010000000000001000000,
31'b1000000000000000000000010000101,
31'b1001001000000000001010000000000,
31'b1010000000000000000010000000000,
31'b1010000000000010000010000000000,
31'b1010000000000100000010000000000,
31'b1010000000000110000010000000000,
31'b0000000010000000000100000000100,
31'b0110000001000000000000001000000,
31'b0010000000000000000000000010011,
31'b0110000001000100000000001000000,
31'b1010000000110000000010000000000,
31'b1001000000000000010000000000001,
31'b0101000000000000010001000001000,
31'b0001000100000000101000000000000,
31'b0010100000100000000000010100000,
31'b1110001000000000000000010000000,
31'b1100010000000000010010000000000,
31'b0001000100001000101000000000000,
31'b1010000000100000000010000000000,
31'b1010000000100010000010000000000,
31'b1101000000000000001000010000000,
31'b0001000100010000101000000000000,
31'b0010001100000000100000000000000,
31'b0110000001100000000000001000000,
31'b0010001100000100100000000000000,
31'b0000000111000000000000000010000,
31'b0000000001000000000000000100011,
31'b0000000000010001010000000000000,
31'b0100000000000010000000001110000,
31'b0100000000000000000000001110000,
31'b0000010000000010000001000100000,
31'b0000010000000000000001000100000,
31'b1000010000100000000000100000100,
31'b0000010000000100000001000100000,
31'b0000000000000011010000000000000,
31'b0000000000000001010000000000000,
31'b0000100001000000000000010010000,
31'b0000000000000101010000000000000,
31'b0000000001000000000100000000100,
31'b0000000000001001010000000000000,
31'b0000000100100010000000000010000,
31'b0000000100100000000000000010000,
31'b0011000000000001000010000000001,
31'b0010000110000000000000000100000,
31'b1000101000000000000000001010000,
31'b0000010010000000010000001000000,
31'b1000010000000100000000100000100,
31'b0000010000100000000001000100000,
31'b1000010000000000000000100000100,
31'b0000000100010000000000000010000,
31'b0001000101000000000000000001000,
31'b0000000000100001010000000000000,
31'b0000100000000000010000000001100,
31'b0000000100001000000000000010000,
31'b0000000100000110000000000010000,
31'b0000000100000100000000000010000,
31'b0000000100000010000000000010000,
31'b0000000100000000000000000010000,
31'b0000000000000000000000000100011,
31'b0000000001010001010000000000000,
31'b0000100000010000000000010010000,
31'b0100100000000001000000100000010,
31'b0000000000010000000100000000100,
31'b0000010001000000000001000100000,
31'b1000000000000000000010000110000,
31'b1000000100000000001001000000100,
31'b0000000000001000000100000000100,
31'b0000000001000001010000000000000,
31'b0000100000000000000000010010000,
31'b0000100000000010000000010010000,
31'b0000000000000000000100000000100,
31'b0000000000000010000100000000100,
31'b0000000000000100000100000000100,
31'b0000000101100000000000000010000,
31'b0001000100010000000000000001000,
31'b1010000000000001000000000001010,
31'b0001000100010100000000000001000,
31'b0001000110000000101000000000000,
31'b0000000100000000001000100100000,
31'b0000010001100000000001000100000,
31'b1000010001000000000000100000100,
31'b0000010000000000001110000000000,
31'b0001000100000000000000000001000,
31'b0001000100000010000000000001000,
31'b0001000100000100000000000001000,
31'b0001000000000000010100010000000,
31'b0000000000100000000100000000100,
31'b0000000101000100000000000010000,
31'b0000000101000010000000000010000,
31'b0000000101000000000000000010000,
31'b1110110000000000000000000000000,
31'b0011100000000000000000000010010,
31'b0100000001000000110000000000000,
31'b0100011000000001000001000000000,
31'b0001000100000000001001000010000,
31'b0001000000000000000010000100100,
31'b1010000000000000100100100000000,
31'b1001000000010000000100000010000,
31'b1000000001000000000100000001000,
31'b1001100000000000000000010000100,
31'b1000100000101000010000000000000,
31'b1001000000001000000100000010000,
31'b1000100000100100010000000000000,
31'b1001000000000100000100000010000,
31'b1000100000100000010000000000000,
31'b1001000000000000000100000010000,
31'b0010000000000000010100000000010,
31'b0010011000000000000000000100000,
31'b0000010000000000000000100001000,
31'b0000010000000010000000100001000,
31'b1100000001000000000000100000010,
31'b0010011000001000000000000100000,
31'b1000100000010000010000000000000,
31'b1000100000010010010000000000000,
31'b1000100000001100010000000000000,
31'b0100001010000000000001001000000,
31'b1000100000001000010000000000000,
31'b1000100000001010010000000000000,
31'b1000100000000100010000000000000,
31'b1000100000000110010000000000000,
31'b1000100000000000010000000000000,
31'b1000100000000010010000000000000,
31'b1000000000010000000100000001000,
31'b1100000010000000000001010000000,
31'b0100000000000000110000000000000,
31'b0100000000000010110000000000000,
31'b1100000000100000000000100000010,
31'b0010110000000000000010001000000,
31'b0100000000001000110000000000000,
31'b0100000000001010110000000000000,
31'b1000000000000000000100000001000,
31'b1000000000000010000100000001000,
31'b1000000000000100000100000001000,
31'b1000000100000000010000010000000,
31'b1000000000001000000100000001000,
31'b1000000000100001000000010010000,
31'b1000100001100000010000000000000,
31'b1001000001000000000100000010000,
31'b1100000000001000000000100000010,
31'b0010011001000000000000000100000,
31'b0100000000100000110000000000000,
31'b0101000000000000000001101000000,
31'b1100000000000000000000100000010,
31'b0010000000000001000000000000110,
31'b1100000000000100000000100000010,
31'b0010010010000000001000000001000,
31'b1000000000100000000100000001000,
31'b1000000000100010000100000001000,
31'b1000100001001000010000000000000,
31'b1000100000000001000100000000100,
31'b0010010000000000100000000000000,
31'b1000000000000001000000010010000,
31'b1000100001000000010000000000000,
31'b1000100001000010010000000000000,
31'b0000000101010000100001000000000,
31'b1100000001000000000001010000000,
31'b0000000001000000000000010001001,
31'b1001000000000000000010010000010,
31'b0000000100000001000000000000101,
31'b0001000000000000000000010010001,
31'b0010000100000000000001100001000,
31'b0001100000010000000000000100010,
31'b0000000101000000100001000000000,
31'b0100001000100000000001001000000,
31'b0010000100000001000010010000000,
31'b0011000000000000000010000010100,
31'b0010000001000000000010000001100,
31'b0001100000000100000000000100010,
31'b1000100010100000010000000000000,
31'b0001100000000000000000000100010,
31'b0011010000000000001000000010000,
31'b1110000000000000001000000000010,
31'b0000010010000000000000100001000,
31'b0000100100001000000000000001001,
31'b1100100100000000000001000000000,
31'b0001010000000000100000000101000,
31'b1000100010010000010000000000000,
31'b0000100100000000000000000001001,
31'b0101000100000001001000000000000,
31'b0100001000000000000001001000000,
31'b1000100010001000010000000000000,
31'b0000100000000000000000101000100,
31'b1000100010000100010000000000000,
31'b0000100000000000100001010000000,
31'b1000100010000000010000000000000,
31'b0000011000000000000000000010000,
31'b0000000100010000100001000000000,
31'b1100000000000000000001010000000,
31'b0000000000000000000000010001001,
31'b1000000000000000101100000000000,
31'b0010000000010000000010000001100,
31'b1100000000001000000001010000000,
31'b0010000000000001100000001000000,
31'b1000010000000000000000011010000,
31'b0000000100000000100001000000000,
31'b0100000000000000011000000001000,
31'b0000000100000100100001000000000,
31'b1000000110000000010000010000000,
31'b0010000000000000000010000001100,
31'b0100100000000000000011000100000,
31'b0010000000010001100000001000000,
31'b0010100000100001000010000000000,
31'b0001100100000000000000000010001,
31'b1100000000100000000001010000000,
31'b0000010000000000100000000110000,
31'b1010000000000001000000010100000,
31'b1100000010000000000000100000010,
31'b0010010000000100001000000001000,
31'b0010010000000010001000000001000,
31'b0010010000000000001000000001000,
31'b0001011000000000000000000001000,
31'b0100001001000000000001001000000,
31'b0001011000000100000000000001000,
31'b0011010000000000000000100100000,
31'b1000001000000000000011000000000,
31'b1000001000000010000011000000000,
31'b1000100011000000010000000000000,
31'b0010100000000001000010000000000,
31'b1100000001000000001000000000001,
31'b0000001010001000000001000100000,
31'b0101010000000000001000001000000,
31'b0000001000100000010000001000000,
31'b0001000000000000001001000010000,
31'b0000001010000000000001000100000,
31'b0010000010000000000001100001000,
31'b0000100010100000000000000001001,
31'b1000100000000001000000000010000,
31'b1000100000000011000000000010000,
31'b1000100000000101000000000010000,
31'b1000000001000000010000010000000,
31'b1001000001100000000000000000100,
31'b0110011000000000000000001000000,
31'b1000100100100000010000000000000,
31'b1001000100000000000100000010000,
31'b0010010000000000000010011000000,
31'b0000001000000100010000001000000,
31'b0000010100000000000000100001000,
31'b0000001000000000010000001000000,
31'b1100100010000000000001000000000,
31'b0000100010000100000000000001001,
31'b1000100100010000010000000000000,
31'b0000100010000000000000000001001,
31'b1001000001001000000000000000100,
31'b1001000000000001010100000000000,
31'b1000100100001000010000000000000,
31'b1000000000000000000000000011100,
31'b1001000001000000000000000000100,
31'b1001000001000010000000000000100,
31'b1000100100000000010000000000000,
31'b1000100100000010010000000000000,
31'b1100000000000000001000000000001,
31'b0000000010000000010100000000001,
31'b0100000100000000110000000000000,
31'b0000000000000000001001000001000,
31'b1100000000001000001000000000001,
31'b0000101000000000000100001001000,
31'b0100000100001000110000000000000,
31'b0000100000000000010010000100000,
31'b0000000010000000100001000000000,
31'b1000000000000100010000010000000,
31'b1000000000000010010000010000000,
31'b1000000000000000010000010000000,
31'b1001000000100000000000000000100,
31'b1001000000100010000000000000100,
31'b1001000000100100000000000000100,
31'b1000000000001000010000010000000,
31'b1100000000100000001000000000001,
31'b0000101000000000001000000100001,
31'b0100001000000001001000100000000,
31'b0000001001000000010000001000000,
31'b1001000000010000000000000000100,
31'b1110010000000000000000010000000,
31'b1100001000000000010010000000000,
31'b0000100011000000000000000001001,
31'b1001000000001000000000000000100,
31'b1001000000001010000000000000100,
31'b1001000000001100000000000000100,
31'b1000000000100000010000010000000,
31'b1001000000000000000000000000100,
31'b1001000000000010000000000000100,
31'b1001000000000100000000000000100,
31'b1001000000000110000000000000100,
31'b0000000001010000100001000000000,
31'b0000001000001000000001000100000,
31'b0010000000010001000010010000000,
31'b0000100000101000000000000001001,
31'b0000000000000001000000000000101,
31'b0000001000000000000001000100000,
31'b0010000000000000000001100001000,
31'b0000100000100000000000000001001,
31'b0000000001000000100001000000000,
31'b0000011000000001010000000000000,
31'b0010000000000001000010010000000,
31'b1000010000000000100010000010000,
31'b0000000001001000100001000000000,
31'b0000010000000000100000000000011,
31'b0010000000010000000001100001000,
31'b0001100100000000000000000100010,
31'b1100100000001000000001000000000,
31'b0000100001000000000011001000000,
31'b1000110000000000000000001010000,
31'b0000100000001000000000000001001,
31'b1100100000000000000001000000000,
31'b0000100000000100000000000001001,
31'b1000001000000000000000100000100,
31'b0000100000000000000000000001001,
31'b0101000000000001001000000000000,
31'b0101000000000011001000000000000,
31'b0110000000000000000101000000010,
31'b1000010000000000010000100000001,
31'b1100100000010000000001000000000,
31'b0000100100000000100001010000000,
31'b1000100110000000010000000000000,
31'b0000100000010000000000000001001,
31'b0000000000010000100001000000000,
31'b0000000000000000010100000000001,
31'b0000000100000000000000010001001,
31'b0000000010000000001001000001000,
31'b0000000001000001000000000000101,
31'b0000001001000000000001000100000,
31'b0010000100000001100000001000000,
31'b0000100010000000010010000100000,
31'b0000000000000000100001000000000,
31'b0000000000000010100001000000000,
31'b0000000000000100100001000000000,
31'b1000000010000000010000010000000,
31'b0000000000001000100001000000000,
31'b0000000000001010100001000000000,
31'b0000000000001100100001000000000,
31'b1001000000000000100000001000010,
31'b0001100000000000000000000010001,
31'b0000100000000000000011001000000,
31'b0001100000000100000000000010001,
31'b0000100001001000000000000001001,
31'b1100100001000000000001000000000,
31'b0000100001000100000000000001001,
31'b1001100000000000000010000000010,
31'b0000100001000000000000000001001,
31'b0000000000100000100001000000000,
31'b0001000000000000010000101000000,
31'b0001000000000000000000010100010,
31'b1000000010100000010000010000000,
31'b1001000010000000000000000000100,
31'b1001000010000010000000000000100,
31'b1001000010000100000000000000100,
31'b0110010000000000000100000000001,
31'b1010000000000000001100000010000,
31'b0010010000100000000000000100000,
31'b0100010000000011000001000000000,
31'b0100010000000001000001000000000,
31'b0000000000000011000000001010000,
31'b0000000000000001000000001010000,
31'b0100000001000001000000000000011,
31'b0100000000010000010000000100000,
31'b1000100000000000001010000000001,
31'b0100000010100000000001001000000,
31'b0100000000001010010000000100000,
31'b0100000000001000010000000100000,
31'b0100000000000110010000000100000,
31'b0100000000000100010000000100000,
31'b0100000000000010010000000100000,
31'b0100000000000000010000000100000,
31'b0010010000000010000000000100000,
31'b0010010000000000000000000100000,
31'b0000011000000000000000100001000,
31'b0000000100000000010000001000000,
31'b0010010000001010000000000100000,
31'b0010010000001000000000000100000,
31'b1000101000010000010000000000000,
31'b0000010010010000000000000010000,
31'b0101000000000000000000010100100,
31'b0100000010000000000001001000000,
31'b1000101000001000010000000000000,
31'b0000010010001000000000000010000,
31'b1000101000000100010000000000000,
31'b0010000000000001010001000000000,
31'b1000101000000000010000000000000,
31'b0000010010000000000000000010000,
31'b1100000000000001000010000010000,
31'b0010010001100000000000000100000,
31'b0100001000000000110000000000000,
31'b0100010001000001000001000000000,
31'b0100000000000101000000000000011,
31'b0000100000000000000000100100010,
31'b0100000000000001000000000000011,
31'b0100000001010000010000000100000,
31'b1000001000000000000100000001000,
31'b1000001000000010000100000001000,
31'b1000001000000100000100000001000,
31'b1010000000000000000100100100000,
31'b1000001000001000000100000001000,
31'b0100100000000000001000001000001,
31'b0100000001000010010000000100000,
31'b0100000001000000010000000100000,
31'b0010010001000010000000000100000,
31'b0010010001000000000000000100000,
31'b0100001000100000110000000000000,
31'b0001010000000000101000000000000,
31'b1100001000000000000000100000010,
31'b0010010001001000000000000100000,
31'b1100000100000000010010000000000,
31'b0001010000001000101000000000000,
31'b0010000000000000000101000000100,
31'b0100100000000000000100000101000,
31'b0010010000000000001000100010000,
31'b0001010000010000101000000000000,
31'b1000000010000000000011000000000,
31'b1000001000000001000000010010000,
31'b1000101001000000010000000000000,
31'b0000010011000000000000000010000,
31'b0110000000000010010000000010000,
31'b0110000000000000010000000010000,
31'b1001000000000000000100100001000,
31'b0110000000000100010000000010000,
31'b0000000100000010000001000100000,
31'b0000000100000000000001000100000,
31'b1000000100100000000000100000100,
31'b0000010000110000000000000010000,
31'b0101000000000000110000100000000,
31'b0100000000100000000001001000000,
31'b1000000000100000000000001001001,
31'b0010000000000001000000001100000,
31'b1000000001100000000011000000000,
31'b0000010000100100000000000010000,
31'b1000000000000000001100000100000,
31'b0000010000100000000000000010000,
31'b0111100000000000000100000000000,
31'b0100000000010000000001001000000,
31'b1000000100001000000000100000100,
31'b0000010000011000000000000010000,
31'b1000000100000100000000100000100,
31'b0000010000010100000000000010000,
31'b1000000100000000000000100000100,
31'b0000010000010000000000000010000,
31'b0100000000000010000001001000000,
31'b0100000000000000000001001000000,
31'b1000000000000000000000001001001,
31'b0000010000001000000000000010000,
31'b1000000001000000000011000000000,
31'b0000010000000100000000000010000,
31'b0000010000000010000000000010000,
31'b0000010000000000000000000010000,
31'b0001100000000100100000000000010,
31'b1100001000000000000001010000000,
31'b0001100000000000100000000000010,
31'b1000100000000000000000110000100,
31'b1000000000110000000011000000000,
31'b1000000000000000000100100010000,
31'b0111000000000000010000000001000,
31'b1000010000000000001001000000100,
31'b0001010000100000000000000001000,
31'b0100001000000000011000000001000,
31'b0001100000010000100000000000010,
31'b0010100000000000000000100010010,
31'b1000000000100000000011000000000,
31'b1000000000100010000011000000000,
31'b1000000001000000001100000100000,
31'b0000010001100000000000000010000,
31'b0001010000010000000000000001000,
31'b0110000000000000000000010001100,
31'b0001100000100000100000000000010,
31'b0001010010000000101000000000000,
31'b1000000000010000000011000000000,
31'b1000000000100000000100100010000,
31'b1000000101000000000000100000100,
31'b0000010001010000000000000010000,
31'b0001010000000000000000000001000,
31'b0100000001000000000001001000000,
31'b0001010000000100000000000001000,
31'b0001000000000000000010001000010,
31'b1000000000000000000011000000000,
31'b1000000000000010000011000000000,
31'b1000000000000100000011000000000,
31'b0000010001000000000000000010000,
31'b0001000000001000000000011000100,
31'b0000000010001000000001000100000,
31'b0001000000000000100001100000000,
31'b0000000000100000010000001000000,
31'b0001000000000000000000011000100,
31'b0000000010000000000001000100000,
31'b1000000010100000000000100000100,
31'b0000000010000100000001000100000,
31'b1010010001000000000010000000000,
31'b0010000000000100000001000010000,
31'b0010000000000010000001000010000,
31'b0010000000000000000001000010000,
31'b0110010000000010000000001000000,
31'b0110010000000000000000001000000,
31'b0110000000000000000010000001010,
31'b0100000100000000010000000100000,
31'b0000000000000110010000001000000,
31'b0000000000000100010000001000000,
31'b0000000000000010010000001000000,
31'b0000000000000000010000001000000,
31'b1001000000000000010001000000010,
31'b0000000010100000000001000100000,
31'b1000000010000000000000100000100,
31'b0000000000001000010000001000000,
31'b0100000000000011000000000110000,
31'b0100000000000001000000000110000,
31'b0000100000000000000000100010001,
31'b0000000000010000010000001000000,
31'b1001001001000000000000000000100,
31'b0110010000100000000000001000000,
31'b1000101100000000010000000000000,
31'b0000010110000000000000000010000,
31'b1100001000000000001000000000001,
31'b0000100000100000001000000100001,
31'b0100001100000000110000000000000,
31'b0000001000000000001001000001000,
31'b0011000000010000000001000001000,
31'b0000100000000000000100001001000,
31'b1100000000100000010010000000000,
31'b0000101000000000010010000100000,
31'b1010010000000000000010000000000,
31'b1010010000000010000010000000000,
31'b1010010000000100000010000000000,
31'b1000001000000000010000010000000,
31'b0011000000000000000001000001000,
31'b0110010001000000000000001000000,
31'b0011000000000100000001000001000,
31'b1111000000000000000000000000001,
31'b0100000000000101001000100000000,
31'b0000100000000000001000000100001,
31'b0100000000000001001000100000000,
31'b0000000001000000010000001000000,
31'b1100000000000100010010000000000,
31'b0000100000100000000100001001000,
31'b1100000000000000010010000000000,
31'b0000000010000000001110000000000,
31'b1010010000100000000010000000000,
31'b0100100000000000000000101000010,
31'b0100100000000000010000010100000,
31'b0000000001010000010000001000000,
31'b1001001000000000000000000000100,
31'b1001001000000010000000000000100,
31'b1100000000010000010010000000000,
31'b0000010111000000000000000010000,
31'b0000000000001010000001000100000,
31'b0000000000001000000001000100000,
31'b1001000000000000000000001100010,
31'b0000000010100000010000001000000,
31'b0000000000000010000001000100000,
31'b0000000000000000000001000100000,
31'b1000000000100000000000100000100,
31'b0000000000000100000001000100000,
31'b0000010000000011010000000000000,
31'b0000010000000001010000000000000,
31'b0010001000000001000010010000000,
31'b0010000010000000000001000010000,
31'b0000010001000000000100000000100,
31'b0000000000010000000001000100000,
31'b1000000100000000001100000100000,
31'b0000010100100000000000000010000,
31'b1000000000001100000000100000100,
31'b0000000010000100010000001000000,
31'b1000000000001000000000100000100,
31'b0000000010000000010000001000000,
31'b1000000000000100000000100000100,
31'b0000000000100000000001000100000,
31'b1000000000000000000000100000100,
31'b0110000000000001000000000000000,
31'b0101001000000001001000000000000,
31'b0100000100000000000001001000000,
31'b1000000100000000000000001001001,
31'b0000010100001000000000000010000,
31'b1000000101000000000011000000000,
31'b0000010100000100000000000010000,
31'b1000000000010000000000100000100,
31'b0000010100000000000000000010000,
31'b0000010000000000000000000100011,
31'b0000001000000000010100000000001,
31'b0001100100000000100000000000010,
31'b0000001010000000001001000001000,
31'b0000010000010000000100000000100,
31'b0000000001000000000001000100000,
31'b1000010000000000000010000110000,
31'b0000000001000100000001000100000,
31'b0000001000000000100001000000000,
31'b0000010001000001010000000000000,
31'b0000110000000000000000010010000,
31'b1010100000000001100000000000000,
31'b0000010000000000000100000000100,
31'b0000010000000010000100000000100,
31'b0000010000000100000100000000100,
31'b0000010101100000000000000010000,
31'b0001101000000000000000000010001,
31'b0000101000000000000011001000000,
31'b1010000000000001000010001000000,
31'b0000000011000000010000001000000,
31'b1000000100010000000011000000000,
31'b0000000001100000000001000100000,
31'b1000000001000000000000100000100,
31'b0000000000000000001110000000000,
31'b0001010100000000000000000001000,
31'b0100000101000000000001001000000,
31'b0001010100000100000000000001000,
31'b0001010000000000010100010000000,
31'b1000000100000000000011000000000,
31'b1000000100000010000011000000000,
31'b1000000100000100000011000000000,
31'b0000010101000000000000000010000,
31'b1111000000000000000000000000000,
31'b0010010000000000000000000010010,
31'b1111000000000100000000000000000,
31'b0011000000000000000001000001001,
31'b1111000000001000000000000000000,
31'b0011000001000000000010001000000,
31'b0000100100000000000100100000100,
31'b1100001000010000001000000000000,
31'b1111000000010000000000000000000,
31'b1000010000000000000000010000100,
31'b0000100000101000001000000100000,
31'b1100001000001000001000000000000,
31'b0000100001000000000111000000000,
31'b1100001000000100001000000000000,
31'b0000100000100000001000000100000,
31'b1100001000000000001000000000000,
31'b1111000000100000000000000000000,
31'b0011101000000000000000000100000,
31'b1000000000000000001010010000000,
31'b1001001000000000000000000000101,
31'b0000100001000010000000100010000,
31'b0000100001000000000000100010000,
31'b0000100000010000001000000100000,
31'b0100000001000000001000011000000,
31'b0000101011000000000000000001000,
31'b1100000000000000010010000000001,
31'b0000100000001000001000000100000,
31'b0100000100000000101010000000000,
31'b0000100000000100001000000100000,
31'b0100000000000100010000000010010,
31'b0000100000000000001000000100000,
31'b0100000000000000010000000010010,
31'b1111000001000000000000000000000,
31'b0011000000001000000010001000000,
31'b1100000000000000101000000100000,
31'b0000101000100000101000000000000,
31'b0010000000000000000001000010001,
31'b0011000000000000000010001000000,
31'b0011010000000000000000000001010,
31'b1110000000000000000000000011000,
31'b0000101010100000000000000001000,
31'b1100000010000000000000000101000,
31'b0000001000000000001010001000000,
31'b0000001010000001000000000000100,
31'b0000100000000000000111000000000,
31'b0011000000010000000010001000000,
31'b0000100001100000001000000100000,
31'b1100001001000000001000000000000,
31'b0000101010010000000000000001000,
31'b0000100000001000000000100010000,
31'b1001000000000000100100000000010,
31'b0000101000000000101000000000000,
31'b0000100000000010000000100010000,
31'b0000100000000000000000100010000,
31'b0100000000000010001000011000000,
31'b0100000000000000001000011000000,
31'b0000101010000000000000000001000,
31'b1000010000000000010000000011000,
31'b0000101010000100000000000001000,
31'b0010100010000000000000100100000,
31'b0000000000000000010000001000001,
31'b0000100000010000000000100010000,
31'b0000100001000000001000000100000,
31'b0100000001000000010000000010010,
31'b1111000010000000000000000000000,
31'b0011000000000000011100000000000,
31'b0000011001000000100000000000010,
31'b0000010000000000000100000000101,
31'b1100001000000000100000000001000,
31'b0000110000000000000000010010001,
31'b0000001000010000010100000000000,
31'b0000010000010000000000000100010,
31'b0000101001100000000000000001000,
31'b1100000001000000000000000101000,
31'b0000001000001000010100000000000,
31'b0000010000001000000000000100010,
31'b0000001000000100010100000000000,
31'b0000010000000100000000000100010,
31'b0000001000000000010100000000000,
31'b0000010000000000000000000100010,
31'b0100000100000000000010000001000,
31'b0110000000000000010000000100010,
31'b1001000100000000000000001010000,
31'b1000000100000000000011000000001,
31'b0110000000000000100001000000100,
31'b0000100000000000100000000101000,
31'b0010101000000000100000100000000,
31'b0001101000010000000000000010000,
31'b0000101001000000000000000001000,
31'b1000000001000000000000100000101,
31'b0000101001000100000000000001000,
31'b0010100001000000000000100100000,
31'b0000101001001000000000000001000,
31'b0001101000000100000000000010000,
31'b0000100010000000001000000100000,
31'b0001101000000000000000000010000,
31'b0000101000110000000000000001000,
31'b1100000000010000000000000101000,
31'b0000011000000000100000000000010,
31'b0000001000010001000000000000100,
31'b0011000000000001001000000000100,
31'b1101000000000000001000100000000,
31'b0000010000000001010000000000001,
31'b0000010001010000000000000100010,
31'b0000101000100000000000000001000,
31'b1100000000000000000000000101000,
31'b0000000000000000000001000100001,
31'b0000001000000001000000000000100,
31'b0000101000101000000000000001000,
31'b1100000000001000000000000101000,
31'b0000001001000000010100000000000,
31'b0000010001000000000000000100010,
31'b0000101000010000000000000001000,
31'b1000000100001000000000001001000,
31'b0001100000000000100000000110000,
31'b0010100000010000000000100100000,
31'b1000011000000000010000100000000,
31'b1000000100000000000000001001000,
31'b1000010100000000000010000000010,
31'b1010000000000000000010110000000,
31'b0000101000000000000000000001000,
31'b1000000000000000000000100000101,
31'b0000101000000100000000000001000,
31'b0010100000000000000000100100000,
31'b0000101000001000000000000001000,
31'b1000000100010000000000001001000,
31'b0000101000001100000000000001000,
31'b0011010000000001000010000000000,
31'b0000000000000000000000110010000,
31'b0100000000010001000000000000010,
31'b0100100000000000001000001000000,
31'b0100100000000010001000001000000,
31'b0100001000000000000101000000000,
31'b0100001000000010000101000000000,
31'b0000100000000000000100100000100,
31'b1000100001000000001010000000000,
31'b0100000000000011000000000000010,
31'b0100000000000001000000000000010,
31'b0100100000010000001000001000000,
31'b0100000000000101000000000000010,
31'b0100001000010000000101000000000,
31'b0100000000001001000000000000010,
31'b0010000010000000000000110100000,
31'b1100001100000000001000000000000,
31'b0100000010000000000010000001000,
31'b0100000010000010000010000001000,
31'b1001000010000000000000001010000,
31'b1000001000000000001000001100000,
31'b0100001000100000000101000000000,
31'b0000000010000000000001000010010,
31'b0010001000000001000100000100000,
31'b0010010000000001010000000000010,
31'b0100000010010000000010000001000,
31'b0100000000100001000000000000010,
31'b0100100000000000000000000001110,
31'b0100000000000000101010000000000,
31'b1011000000000000000000001100000,
31'b0100001000000000000010100010000,
31'b0010000000000000110000000000100,
31'b0100000100000000010000000010010,
31'b0100000000000000010000000100001,
31'b0100000001010001000000000000010,
31'b0100100001000000001000001000000,
31'b0000100000000001010000100000000,
31'b0100001001000000000101000000000,
31'b1000100000000100001010000000000,
31'b1000100000000010001010000000000,
31'b1000100000000000001010000000000,
31'b0100000001000011000000000000010,
31'b0100000001000001000000000000010,
31'b0000000000000010001000010100000,
31'b0000000000000000001000010100000,
31'b1000110000100000000000000000100,
31'b1000010000000101000000000001000,
31'b1000010000000011000000000001000,
31'b1000010000000001000000000001000,
31'b0000010010000000000000000010001,
31'b1000101000000000010000000000001,
31'b0010010000000000000100000000110,
31'b0010001000000000010000000100100,
31'b1000110000010000000000000000100,
31'b1000000010000000000000001001000,
31'b1000010010000000000010000000010,
31'b1000100000100000001010000000000,
31'b1000110000001000000000000000100,
31'b0111000000000000000010000100000,
31'b1000010000000000000100010010000,
31'b0010000000000001100100000000000,
31'b1000110000000000000000000000100,
31'b1000110000000010000000000000100,
31'b1000000000000000101000001000000,
31'b1000010000100001000000000001000,
31'b0100000000100000000010000001000,
31'b0100000010010001000000000000010,
31'b1010100000000000000010100000000,
31'b1000100000000000010100001000000,
31'b0100001010000000000101000000000,
31'b0000001000010000000000010001000,
31'b0010100000000001011000000000000,
31'b0001010000100000000000000001001,
31'b0100000010000011000000000000010,
31'b0100000010000001000000000000010,
31'b1011000000000000010001000000000,
31'b0100010000000000001000000001100,
31'b0000001000000010000000010001000,
31'b0000001000000000000000010001000,
31'b0010000000000000000000110100000,
31'b0000010100000000000000000100010,
31'b0100000000000000000010000001000,
31'b0100000000000010000010000001000,
31'b1001000000000000000000001010000,
31'b1000000000000000000011000000001,
31'b0100000000001000000010000001000,
31'b0000000000000000000001000010010,
31'b1001000000001000000000001010000,
31'b0001010000000000000000000001001,
31'b0100000000010000000010000001000,
31'b0100000010100001000000000000010,
31'b1001000000010000000000001010000,
31'b1010000000000000100000101000000,
31'b0100000000011000000010000001000,
31'b0000001000100000000000010001000,
31'b0010000010000000110000000000100,
31'b0001101100000000000000000010000,
31'b0000010000100000000000000010001,
31'b1000000000101000000000001001000,
31'b0001001000010000000000010010000,
31'b0010100000000000001100000000100,
31'b1000010000000001101000000000000,
31'b1000000000100000000000001001000,
31'b1000100000000001000000001000100,
31'b1000100010000000001010000000000,
31'b0001110000000000100001000000000,
31'b1100000100000000000000000101000,
31'b0001001000000000000000010010000,
31'b0000001100000001000000000000100,
31'b1000100000000000100010000001000,
31'b1000000000000000001000000000110,
31'b0110000000000000010000000010001,
31'b1000010010000001000000000001000,
31'b0000010000000000000000000010001,
31'b1000000000001000000000001001000,
31'b0001000000000000000001000001010,
31'b1000000001000000000011000000001,
31'b1000000000000010000000001001000,
31'b1000000000000000000000001001000,
31'b1000010000000000000010000000010,
31'b1000000000000100000000001001000,
31'b0000101100000000000000000001000,
31'b1000000100000000000000100000101,
31'b0001001000100000000000010010000,
31'b0010100100000000000000100100000,
31'b1000110010000000000000000000100,
31'b1000000000010000000000001001000,
31'b1000010000010000000010000000010,
31'b1000000000010100000000001001000,
31'b1111001000000000000000000000000,
31'b0011100000100000000000000100000,
31'b0000010100000000000100001010000,
31'b1100000000011000001000000000000,
31'b1000000000000000010000010000001,
31'b1100000000010100001000000000000,
31'b0000000100000000101000010000000,
31'b1100000000010000001000000000000,
31'b0000100011100000000000000001000,
31'b1100000000001100001000000000000,
31'b0000000010001000010100000000000,
31'b1100000000001000001000000000000,
31'b0000000010000100010100000000000,
31'b1100000000000100001000000000000,
31'b0000000010000000010100000000000,
31'b1100000000000000001000000000000,
31'b0110010010000000000100000000000,
31'b0011100000000000000000000100000,
31'b1001000000000010000000000000101,
31'b1001000000000000000000000000101,
31'b1100010000000000000010000000100,
31'b0011100000001000000000000100000,
31'b0010100010000000100000100000000,
31'b1100000000110000001000000000000,
31'b0000100011000000000000000001000,
31'b0011100000010000000000000100000,
31'b0000101000001000001000000100000,
31'b1100000000101000001000000000000,
31'b0000101000000100001000000100000,
31'b1100000000100100001000000000000,
31'b0000101000000000001000000100000,
31'b1100000000100000001000000000000,
31'b0000100010110000000000000001000,
31'b0000100000000001000010000000010,
31'b0000010010000000100000000000010,
31'b0000100000100000101000000000000,
31'b1100000000000000000000100110000,
31'b0011001000000000000010001000000,
31'b0001010000000000010000011000000,
31'b1100000001010000001000000000000,
31'b0000100010100000000000000001000,
31'b0000010000000000001000000001010,
31'b0000000000000000001010001000000,
31'b0000000010000001000000000000100,
31'b0000101000000000000111000000000,
31'b1100000001000100001000000000000,
31'b0000000011000000010100000000000,
31'b1100000001000000001000000000000,
31'b0000100010010000000000000001000,
31'b0000010000000000000000001000100,
31'b0000100000000010101000000000000,
31'b0000100000000000101000000000000,
31'b1000010010000000010000100000000,
31'b0000101000000000000000100010000,
31'b0100000100000000001010000100000,
31'b0100000000000000000001000010100,
31'b0000100010000000000000000001000,
31'b0000100010000010000000000001000,
31'b0000100010000100000000000001000,
31'b0000100000010000101000000000000,
31'b0000100010001000000000000001000,
31'b0000101000010000000000100010000,
31'b0000101001000000001000000100000,
31'b1100000001100000001000000000000,
31'b1100000000001000100000000001000,
31'b0000000100011000000000010001000,
31'b0000010001000000100000000000010,
31'b0000000001010001000000000000100,
31'b1100000000000000100000000001000,
31'b0000000100010000000000010001000,
31'b0000000000010000010100000000000,
31'b0000000000000000100001000000001,
31'b0000100001100000000000000001000,
31'b0000000100001000000000010001000,
31'b0000000000001000010100000000000,
31'b0000000001000001000000000000100,
31'b0000000000000100010100000000000,
31'b0000000100000000000000010001000,
31'b0000000000000000010100000000000,
31'b0000000000000010010100000000000,
31'b0110010000000000000100000000000,
31'b0110010000000010000100000000000,
31'b0110010000000100000100000000000,
31'b1001000010000000000000000000101,
31'b1100000000100000100000000001000,
31'b0001100000010100000000000010000,
31'b0010100000000000100000100000000,
31'b0001100000010000000000000010000,
31'b0000100001000000000000000001000,
31'b0001000000000000000100010000100,
31'b0000100001000100000000000001000,
31'b0001100000001000000000000010000,
31'b0000100001001000000000000001000,
31'b0001100000000100000000000010000,
31'b0000000000100000010100000000000,
31'b0001100000000000000000000010000,
31'b0000100000110000000000000001000,
31'b0000000000010101000000000000100,
31'b0000010000000000100000000000010,
31'b0000000000010001000000000000100,
31'b1100000001000000100000000001000,
31'b0010000100000000000001001000100,
31'b0000010000001000100000000000010,
31'b0000000001000000100001000000001,
31'b0000100000100000000000000001000,
31'b0000000000000101000000000000100,
31'b0000000000000011000000000000100,
31'b0000000000000001000000000000100,
31'b0000100000101000000000000001000,
31'b0000000101000000000000010001000,
31'b0000000001000000010100000000000,
31'b0000000000001001000000000000100,
31'b0000100000010000000000000001000,
31'b0000100000010010000000000001000,
31'b0000100000010100000000000001000,
31'b0000100010000000101000000000000,
31'b1000010000000000010000100000000,
31'b1000010000000010010000100000000,
31'b1010000000000000000100000001010,
31'b0101000000000001001000000000001,
31'b0000100000000000000000000001000,
31'b0000100000000010000000000001000,
31'b0000100000000100000000000001000,
31'b0000000000100001000000000000100,
31'b0000100000001000000000000001000,
31'b0000100000001010000000000001000,
31'b0000100000001100000000000001000,
31'b0001100001000000000000000010000,
31'b0100000000001000000101000000000,
31'b0100001000010001000000000000010,
31'b0000010000000000000100001010000,
31'b1000000000100000001000001100000,
31'b0100000000000000000101000000000,
31'b0100000000000010000101000000000,
31'b0000000000000000101000010000000,
31'b1000000000000000000100000001001,
31'b0100001000000011000000000000010,
31'b0100001000000001000000000000010,
31'b0001010000000000110010000000000,
31'b1100000100001000001000000000000,
31'b0100000000010000000101000000000,
31'b0000000010000000000000010001000,
31'b0000000110000000010100000000000,
31'b1100000100000000001000000000000,
31'b0100001010000000000010000001000,
31'b1000100001000000010000000000001,
31'b1000000000000010001000001100000,
31'b1000000000000000001000001100000,
31'b0100000000100000000101000000000,
31'b0100000000100010000101000000000,
31'b0010000000000001000100000100000,
31'b1000000000100000000100000001001,
31'b0000000010000001000100000010000,
31'b0100001000100001000000000000010,
31'b0010010000000000010101000000000,
31'b1100000000000000000000100000011,
31'b0100000000110000000101000000000,
31'b0100000000000000000010100010000,
31'b0010001000000000110000000000100,
31'b1100000100100000001000000000000,
31'b1010000000000000010001100000000,
31'b1000100000100000010000000000001,
31'b0001000010010000000000010010000,
31'b0010000010000000100000110000000,
31'b0100000001000000000101000000000,
31'b0100010000010000000000000100100,
31'b0001000000000000000110000000010,
31'b1000101000000000001010000000000,
31'b1011100000000000000010000000000,
31'b0100010000001000000000000100100,
31'b0001000010000000000000010010000,
31'b0000001000000000001000010100000,
31'b0100010000000010000000000100100,
31'b0100010000000000000000000100100,
31'b0001000010001000000000010010000,
31'b1100000101000000001000000000000,
31'b1000100000000010010000000000001,
31'b1000100000000000010000000000001,
31'b0100100000000000010001000001000,
31'b0010000000000000010000000100100,
31'b0100000001100000000101000000000,
31'b1000100000001000010000000000001,
31'b0100000000000000001010000100000,
31'b0100000100000000000001000010100,
31'b1000000000000000000000101010000,
31'b1000100000010000010000000000001,
31'b1100100000000000001000010000000,
31'b0010001000000001100100000000000,
31'b1000111000000000000000000000100,
31'b0000010000000000000000100001001,
31'b1100010000000000000001100000000,
31'b0010010000000001000001000000100,
31'b0100001000100000000010000001000,
31'b0000000000011000000000010001000,
31'b0001000001010000000000010010000,
31'b0010000001000000100000110000000,
31'b0100000010000000000101000000000,
31'b0000000000010000000000010001000,
31'b0000000100010000010100000000000,
31'b0000000100000000100001000000001,
31'b0000000000100001000100000010000,
31'b0000000000001000000000010001000,
31'b0001000001000000000000010010000,
31'b0000000101000001000000000000100,
31'b0000000000000010000000010001000,
31'b0000000000000000000000010001000,
31'b0000000100000000010100000000000,
31'b0000000000000100000000010001000,
31'b0100001000000000000010000001000,
31'b0100001000000010000010000001000,
31'b1001001000000000000000001010000,
31'b1000001000000000000011000000001,
31'b0100001000001000000010000001000,
31'b0000001000000000000001000010010,
31'b0010100100000000100000100000000,
31'b0001100100010000000000000010000,
31'b0000000000000001000100000010000,
31'b0000000000101000000000010001000,
31'b0001000000000000010000000001100,
31'b0001100100001000000000000010000,
31'b0000000000100010000000010001000,
31'b0000000000100000000000010001000,
31'b0000100000000001000000010000100,
31'b0001100100000000000000000010000,
31'b0001100000000000000000000100011,
31'b0010000000001000000001001000100,
31'b0001000000010000000000010010000,
31'b0010000000000000100000110000000,
31'b0100100000000000000000001101000,
31'b0010000000000000000001001000100,
31'b0001000010000000000110000000010,
31'b0010000000001000100000110000000,
31'b0001000000000100000000010010000,
31'b0000000100000101000000000000100,
31'b0001000000000000000000010010000,
31'b0000000100000001000000000000100,
31'b0001100000000000000100000000100,
31'b0000000001000000000000010001000,
31'b0001000000001000000000010010000,
31'b0000000100001001000000000000100,
31'b0000100100010000000000000001000,
31'b1000100010000000010000000000001,
31'b0001001000000000000001000001010,
31'b0010000010000000010000000100100,
31'b1000010100000000010000100000000,
31'b1000001000000000000000001001000,
31'b1010000000000000000000101100000,
31'b1000001000000100000000001001000,
31'b0000100100000000000000000001000,
31'b0000100100000010000000000001000,
31'b0001000000100000000000010010000,
31'b0000100000000000010100010000000,
31'b0000100100001000000000000001000,
31'b0000000000000000010000000010100,
31'b0001000000101000000000010010000,
31'b0001000000000001000100000001000,
31'b0100000100000000100000000000100,
31'b0010000000000000000000000010010,
31'b0110000001000000000000001000001,
31'b0010000000000100000000000010010,
31'b0110000000000000000011000001000,
31'b0010000000001000000000000010010,
31'b1010000000000010000010000000001,
31'b1010000000000000000010000000001,
31'b1000000000000010000000010000100,
31'b1000000000000000000000010000100,
31'b1001000000101000010000000000000,
31'b1000000000000100000000010000100,
31'b1001000000100100010000000000000,
31'b1000000000001000000000010000100,
31'b1001000000100000010000000000000,
31'b0000000010000000000000000100010,
31'b0110001010000000000100000000000,
31'b0010000000100000000000000010010,
31'b1001000000011000010000000000000,
31'b0100000110000000000000001000010,
31'b1100001000000000000010000000100,
31'b0010001000000001000010100000000,
31'b1001000000010000010000000000000,
31'b1010000000100000000010000000001,
31'b1001000000001100010000000000000,
31'b1000000000100000000000010000100,
31'b1001000000001000010000000000000,
31'b1001000000001010010000000000000,
31'b1001000000000100010000000000000,
31'b1001000000000110010000000000000,
31'b1001000000000000010000000000000,
31'b1001000000000010010000000000000,
31'b0110000000000100000000001000001,
31'b0010000001000000000000000010010,
31'b0110000000000000000000001000001,
31'b0110000000000010000000001000001,
31'b0011000000000100000000000001010,
31'b0011010000000000000010001000000,
31'b0011000000000000000000000001010,
31'b1010000001000000000010000000001,
31'b1001100000000000000100000001000,
31'b1000000001000000000000010000100,
31'b0110000000010000000000001000001,
31'b1000000100001001000000000001000,
31'b1000100100100000000000000000100,
31'b1000000100000101000000000001000,
31'b1001000001100000010000000000000,
31'b1000000100000001000000000001000,
31'b0000001000000010000000001000100,
31'b0000001000000000000000001000100,
31'b0110000000100000000000001000001,
31'b0100000000000000100100000010000,
31'b1000100100010000000000000000100,
31'b0000110000000000000000100010000,
31'b1001000001010000010000000000000,
31'b0100010000000000001000011000000,
31'b1000100100001000000000000000100,
31'b1000000000000000010000000011000,
31'b1001000001001000010000000000000,
31'b1001000000000001000100000000100,
31'b1000100100000000000000000000100,
31'b1000100100000010000000000000100,
31'b1001000001000000010000000000000,
31'b1001000001000010010000000000000,
31'b0110001000100000000100000000000,
31'b0010000010000000000000000010010,
31'b0000001001000000100000000000010,
31'b0000000000000000000100000000101,
31'b0000100000000010000000010010001,
31'b0000100000000000000000010010001,
31'b0000000001000001010000000000001,
31'b0000000000010000000000000100010,
31'b1001000000000000000001001100000,
31'b1000000010000000000000010000100,
31'b0000000000001010000000000100010,
31'b0000000000001000000000000100010,
31'b0000000000000110000000000100010,
31'b0000000000000100000000000100010,
31'b0000000000000010000000000100010,
31'b0000000000000000000000000100010,
31'b0110001000000000000100000000000,
31'b0110001000000010000100000000000,
31'b0110001000000100000100000000000,
31'b0100000100000000000000001000010,
31'b1101000100000000000001000000000,
31'b0001000100000100000000000001001,
31'b1001000010010000010000000000000,
31'b0001000100000000000000000001001,
31'b0110001000010000000100000000000,
31'b1000000010100000000000010000100,
31'b1001000010001000010000000000000,
31'b0001000000000000000000101000100,
31'b1001000010000100010000000000000,
31'b0001000000000000100001010000000,
31'b1001000010000000010000000000000,
31'b0000000000100000000000000100010,
31'b0000001000000100100000000000010,
31'b0010000100000000100100001000000,
31'b0000001000000000100000000000010,
31'b0000001000000010100000000000010,
31'b0000000000000101010000000000001,
31'b0100100000000000010000100100000,
31'b0000000000000001010000000000001,
31'b0000000001010000000000000100010,
31'b0001100100000000100001000000000,
31'b1100010000000000000000000101000,
31'b0000010000000000000001000100001,
31'b0000011000000001000000000000100,
31'b0100000000000011001000010000000,
31'b0100000000000001001000010000000,
31'b0000000001000010000000000100010,
31'b0000000001000000000000000100010,
31'b0000000100000000000000000010001,
31'b0000001010000000000000001000100,
31'b0000001000100000100000000000010,
31'b0100000101000000000000001000010,
31'b1000001000000000010000100000000,
31'b1000010100000000000000001001000,
31'b1000000100000000000010000000010,
31'b1010000000000000010000000101000,
31'b0000111000000000000000000001000,
31'b1000010000000000000000100000101,
31'b0000111000000100000000000001000,
31'b0011000000001001000010000000000,
31'b1000100110000000000000000000100,
31'b0110000000000000100100000100000,
31'b1001000011000000010000000000000,
31'b0011000000000001000010000000000,
31'b0100000000000000100000000000100,
31'b0100000000000010100000000000100,
31'b0100000000000100100000000000100,
31'b0100000010100000000000001000010,
31'b0100000000001000100000000000100,
31'b0100000000001010100000000000100,
31'b0100000000001100100000000000100,
31'b1010000100000000000010000000001,
31'b1001000000000001000000000010000,
31'b1000000100000000000000010000100,
31'b1001000000000101000000000010000,
31'b1000000100000100000000010000100,
31'b1001000000001001000000000010000,
31'b1000000100001000000000010000100,
31'b1001000100100000010000000000000,
31'b1000000001000001000000000001000,
31'b0100000000100000100000000000100,
31'b0100000010000100000000001000010,
31'b0100000010000010000000001000010,
31'b0100000010000000000000001000010,
31'b1101000010000000000001000000000,
31'b0010000000000101010000000000010,
31'b1001000100010000010000000000000,
31'b0010000000000001010000000000010,
31'b1001000000100001000000000010000,
31'b1000100000000001010100000000000,
31'b1001000100001000010000000000000,
31'b0100010000000000101010000000000,
31'b1000100001000000000000000000100,
31'b1001000000000000000100010001000,
31'b1001000100000000010000000000000,
31'b1001000100000010010000000000000,
31'b0100000001000000100000000000100,
31'b0100001000000000000100000000011,
31'b0110000100000000000000001000001,
31'b1000000000011001000000000001000,
31'b1000100000110000000000000000100,
31'b1000000000010101000000000001000,
31'b1000000010100000000010000000010,
31'b1000000000010001000000000001000,
31'b1001000001000001000000000010000,
31'b1000000101000000000000010000100,
31'b1000000000100000000100010010000,
31'b1000000000001001000000000001000,
31'b1000100000100000000000000000100,
31'b1000000000000101000000000001000,
31'b1000000000000011000000000001000,
31'b1000000000000001000000000001000,
31'b0000000010000000000000000010001,
31'b0000001100000000000000001000100,
31'b0010000000000000000100000000110,
31'b0100000100000000100100000010000,
31'b1000100000010000000000000000100,
31'b1000100000010010000000000000100,
31'b1000000010000000000010000000010,
31'b1000000010000010000010000000010,
31'b1000100000001000000000000000100,
31'b1000100000001010000000000000100,
31'b1000000000000000000100010010000,
31'b1000000000101001000000000001000,
31'b1000100000000000000000000000100,
31'b1000100000000010000000000000100,
31'b0010000000000000000000000100001,
31'b1000000000100001000000000001000,
31'b0100000010000000100000000000100,
31'b0100000010000010100000000000100,
31'b0100000010000100100000000000100,
31'b0100000000100000000000001000010,
31'b1101000000100000000001000000000,
31'b0001101000000000000001000100000,
31'b1011000000000001000000000100000,
31'b0001000000100000000000000001001,
31'b1001000010000001000000000010000,
31'b1000001000000001001000000100000,
31'b0100100000000000100010000000010,
31'b0100000000000000001000000001100,
31'b0010001000000000000100001100000,
31'b0000011000000000000000010001000,
31'b0010000000000000010010000001000,
31'b0000000100000000000000000100010,
31'b0000000001000000000000000010001,
31'b0100000000000100000000001000010,
31'b0100000000000010000000001000010,
31'b0100000000000000000000001000010,
31'b1101000000000000000001000000000,
31'b0001000000000100000000000001001,
31'b1000000001000000000010000000010,
31'b0001000000000000000000000001001,
31'b0100100000000001001000000000000,
31'b0100100000000011001000000000000,
31'b0100100000000101001000000000000,
31'b0100000000010000000000001000010,
31'b1101000000010000000001000000000,
31'b0001000100000000100001010000000,
31'b1001000110000000010000000000000,
31'b0001000000010000000000000001001,
31'b0000000000100000000000000010001,
31'b0010000000000000100100001000000,
31'b0000001100000000100000000000010,
31'b0110001000000000000000000010100,
31'b1000000000000001101000000000000,
31'b1000010000100000000000001001000,
31'b1000000000100000000010000000010,
31'b1000000010010001000000000001000,
31'b0001100000000000100001000000000,
31'b0011000000000000010010000010000,
31'b0001100000000100100001000000000,
31'b1100001000000000000000010000010,
31'b1000100010100000000000000000100,
31'b1000010000000000001000000000110,
31'b1000000010000011000000000001000,
31'b1000000010000001000000000001000,
31'b0000000000000000000000000010001,
31'b0000000000000010000000000010001,
31'b0000000000000100000000000010001,
31'b0100000001000000000000001000010,
31'b0000000000001000000000000010001,
31'b1000010000000000000000001001000,
31'b1000000000000000000010000000010,
31'b1000000000000010000010000000010,
31'b0000000000010000000000000010001,
31'b0000100000000000010000101000000,
31'b0000100000000000000000010100010,
31'b0100000001010000000000001000010,
31'b1000100010000000000000000000100,
31'b1000100010000010000000000000100,
31'b1000000000010000000010000000010,
31'b1000000010100001000000000001000,
31'b0110000010100000000100000000000,
31'b0010001000000000000000000010010,
31'b0000000100000000000100001010000,
31'b0010001000000100000000000010010,
31'b1100000000100000000010000000100,
31'b0010001000001000000000000010010,
31'b0001000001000000010000011000000,
31'b1100010000010000001000000000000,
31'b1001000000000000001010000000001,
31'b1000001000000000000000010000100,
31'b0001000100000000110010000000000,
31'b1100010000001000001000000000000,
31'b0010000010000000000000100001010,
31'b1100010000000100001000000000000,
31'b0001000000000000001000000010010,
31'b1100010000000000001000000000000,
31'b0110000010000000000100000000000,
31'b0000000001000000000000001000100,
31'b0110000010000100000100000000000,
31'b0010000100000000100000000000001,
31'b1100000000000000000010000000100,
31'b0010000000000001000010100000000,
31'b1100000000000100000010000000100,
31'b0010000100001000100000000000001,
31'b0110000010010000000100000000000,
31'b0010000000000000000001010001000,
31'b1110000000000000000000010000001,
31'b0010000100010000100000000000001,
31'b1100000000010000000010000000100,
31'b0010000000010001000010100000000,
31'b1001001000000000010000000000000,
31'b1100010000100000001000000000000,
31'b0000000010000100100000000000010,
31'b0000000000100000000000001000100,
31'b0000000010000000100000000000010,
31'b0000000010000010100000000000010,
31'b1000000010100000010000100000000,
31'b0001000000000000000000100100010,
31'b0001000000000000010000011000000,
31'b0001000000000100000000100100010,
31'b0000100000000000100010000000100,
31'b0000000000000000001000000001010,
31'b0000010000000000001010001000000,
31'b0000010010000001000000000000100,
31'b0100000100000010000000000100100,
31'b0100000100000000000000000100100,
31'b0001000001000000001000000010010,
31'b1100010001000000001000000000000,
31'b0000000000000010000000001000100,
31'b0000000000000000000000001000100,
31'b0000000010100000100000000000010,
31'b0000000000000100000000001000100,
31'b1000000010000000010000100000000,
31'b0000000000001000000000001000100,
31'b1001000000000000000001000000110,
31'b0000000000001100000000001000100,
31'b0000110010000000000000000001000,
31'b0000000000010000000000001000100,
31'b0000110010000100000000000001000,
31'b0000000000010100000000001000100,
31'b1000101100000000000000000000100,
31'b0000000100000000000000100001001,
31'b1100000100000000000001100000000,
31'b0010000100000001000001000000100,
31'b0110000000100000000100000000000,
31'b0110000000100010000100000000000,
31'b0000000001000000100000000000010,
31'b0000001000000000000100000000101,
31'b1100010000000000100000000001000,
31'b0001100100000000000001000100000,
31'b0000010000010000010100000000000,
31'b0000010000000000100001000000001,
31'b0110000000110000000100000000000,
31'b1000001010000000000000010000100,
31'b0000010000001000010100000000000,
31'b0000010001000001000000000000100,
31'b0010000000000000000000100001010,
31'b0000010100000000000000010001000,
31'b0000010000000000010100000000000,
31'b0000001000000000000000000100010,
31'b0110000000000000000100000000000,
31'b0110000000000010000100000000000,
31'b0110000000000100000100000000000,
31'b0110000000000110000100000000000,
31'b1000000001000000010000100000000,
31'b1100000000000001001000001000000,
31'b1100100000010000000000000000010,
31'b0001110000010000000000000010000,
31'b0110000000010000000100000000000,
31'b0110000000010010000100000000000,
31'b1100100000001000000000000000010,
31'b0001110000001000000000000010000,
31'b1100100000000100000000000000010,
31'b0001110000000100000000000010000,
31'b1100100000000000000000000000010,
31'b0001110000000000000000000010000,
31'b0000000000000100100000000000010,
31'b0000000010100000000000001000100,
31'b0000000000000000100000000000010,
31'b0000000000000010100000000000010,
31'b1000000000100000010000100000000,
31'b1001000000000000100001001000000,
31'b0000000000001000100000000000010,
31'b0000000000001010100000000000010,
31'b0000110000100000000000000001000,
31'b0000010000000101000000000000100,
31'b0000000000010000100000000000010,
31'b0000010000000001000000000000100,
31'b1010100000000000100100000000000,
31'b0100001000000001001000010000000,
31'b0000010001000000010100000000000,
31'b0000010000001001000000000000100,
31'b0000000000000001001010000000000,
31'b0000000010000000000000001000100,
31'b0000000000100000100000000000010,
31'b0000000010000100000000001000100,
31'b1000000000000000010000100000000,
31'b1000000000000010010000100000000,
31'b1000000000000100010000100000000,
31'b1000000000000110010000100000000,
31'b0000110000000000000000000001000,
31'b0000110000000010000000000001000,
31'b0000110000000100000000000001000,
31'b0000100000000000000010001000010,
31'b1000000000010000010000100000000,
31'b1000100000000000000000001010001,
31'b1100100001000000000000000000010,
31'b0011001000000001000010000000000,
31'b0100001000000000100000000000100,
31'b0100001000000010100000000000100,
31'b0000000000000000000100001010000,
31'b0010000000100000100000000000001,
31'b0100010000000000000101000000000,
31'b0100010000000010000101000000000,
31'b0000010000000000101000010000000,
31'b1010000000000001001000000010000,
31'b1001001000000001000000000010000,
31'b1000001100000000000000010000100,
31'b0001000000000000110010000000000,
31'b0011100000000000000001000010000,
31'b0100010000010000000101000000000,
31'b0100000001000000000000000100100,
31'b0001000100000000001000000010010,
31'b1100010100000000001000000000000,
31'b0110000110000000000100000000000,
31'b0010000000000100100000000000001,
31'b0010000000000010100000000000001,
31'b0010000000000000100000000000001,
31'b1100000100000000000010000000100,
31'b0010000100000001000010100000000,
31'b0010010000000001000100000100000,
31'b0010000000001000100000000000001,
31'b0010000010000000001000000001001,
31'b0010000100000000000001010001000,
31'b0010000000000000010101000000000,
31'b0010000000010000100000000000001,
31'b1001000000000000000010100000010,
31'b0000000001000000000000100001001,
31'b1100000001000000000001100000000,
31'b0010000001000001000001000000100,
31'b0100001001000000100000000000100,
31'b0100000000000000000100000000011,
31'b0000000110000000100000000000010,
31'b0110000010000000000000000010100,
31'b0100010001000000000101000000000,
31'b0100000000010000000000000100100,
31'b0001010000000000000110000000010,
31'b1100000000000000000110000010000,
31'b0100000000001010000000000100100,
31'b0100000000001000000000000100100,
31'b0001010010000000000000010010000,
31'b1100000010000000000000010000010,
31'b0100000000000010000000000100100,
31'b0100000000000000000000000100100,
31'b1100000000100000000001100000000,
31'b1000001000000001000000000001000,
31'b0000001010000000000000000010001,
31'b0000000100000000000000001000100,
31'b0010001000000000000100000000110,
31'b0010000001000000100000000000001,
31'b1000101000010000000000000000100,
31'b0000000100001000000000001000100,
31'b1100000000010000000001100000000,
31'b0010000001001000100000000000001,
31'b1000101000001000000000000000100,
31'b0000000100010000000000001000100,
31'b1100000000001000000001100000000,
31'b0010000001010000100000000000001,
31'b1000101000000000000000000000100,
31'b0000000000000000000000100001001,
31'b1100000000000000000001100000000,
31'b0010000000000001000001000000100,
31'b0110000100100000000100000000000,
31'b1000100000000000010000110000000,
31'b0000000101000000100000000000010,
31'b0110000001000000000000000010100,
31'b0111000000000000000000000001100,
31'b0001100000000000000001000100000,
31'b0000010100010000010100000000000,
31'b0001100000000100000001000100000,
31'b1000000000000011001000000100000,
31'b1000000000000001001000000100000,
31'b0001010001000000000000010010000,
31'b1100000001000000000000010000010,
31'b0010000000000000000100001100000,
31'b0000010000000000000000010001000,
31'b0000010100000000010100000000000,
31'b0000010000000100000000010001000,
31'b0110000100000000000100000000000,
31'b0110000100000010000100000000000,
31'b0110000100000100000100000000000,
31'b0100001000000000000000001000010,
31'b1101001000000000000001000000000,
31'b0001100000100000000001000100000,
31'b1001100000000000000000100000100,
31'b0001001000000000000000000001001,
31'b0010000000000000001000000001001,
31'b1010000000000000100100010000000,
31'b0010000010000000010101000000000,
31'b1110000000000000001001000000000,
31'b0010000000100000000100001100000,
31'b0000010000100000000000010001000,
31'b1100100100000000000000000000010,
31'b0001110100000000000000000010000,
31'b0000001000100000000000000010001,
31'b0110000000000100000000000010100,
31'b0000000100000000100000000000010,
31'b0110000000000000000000000010100,
31'b1000001000000001101000000000000,
31'b0110100000000000000100010000000,
31'b0000000100001000100000000000010,
31'b0110000000001000000000000010100,
31'b0001101000000000100001000000000,
31'b1100000000000100000000010000010,
31'b0001010000000000000000010010000,
31'b1100000000000000000000010000010,
31'b0101000000000000000001011000000,
31'b0100000010000000000000000100100,
31'b0001010000001000000000010010000,
31'b1100000000001000000000010000010,
31'b0000001000000000000000000010001,
31'b0000001000000010000000000010001,
31'b0000001000000100000000000010001,
31'b0110000000100000000000000010100,
31'b1000000100000000010000100000000,
31'b1000011000000000000000001001000,
31'b1000001000000000000010000000010,
31'b1000001000000010000010000000010,
31'b0000110100000000000000000001000,
31'b0000110100000010000000000001000,
31'b0001010000100000000000010010000,
31'b1100000000100000000000010000010,
31'b1000101010000000000000000000100,
31'b0000010000000000010000000010100,
31'b1100000010000000000001100000000,
31'b0011000000000000001000000010001,
31'b1111100000000000000000000000000,
31'b0011001000100000000000000100000,
31'b0100000100000000001000001000000,
31'b0101001000000001000001000000000,
31'b0000010100000000001001000010000,
31'b0000010000000000000010000100100,
31'b0000000100000000000100100000100,
31'b1000010000010000000100000010000,
31'b0000001011100000000000000001000,
31'b1100000000000000000101001000000,
31'b0000000000101000001000000100000,
31'b1000010000001000000100000010000,
31'b0000000001000000000111000000000,
31'b1000010000000100000100000010000,
31'b0000000000100000001000000100000,
31'b1000010000000000000100000010000,
31'b0010000010000000001000000010000,
31'b0011001000000000000000000100000,
31'b0001000000000000000000100001000,
31'b0001000000000010000000100001000,
31'b0000000001000010000000100010000,
31'b0000000001000000000000100010000,
31'b0000000000010000001000000100000,
31'b0000000001000100000000100010000,
31'b0000001011000000000000000001000,
31'b0011001000010000000000000100000,
31'b0000000000001000001000000100000,
31'b0010000000000000100000000011000,
31'b0000000000000100001000000100000,
31'b0000000001010000000000100010000,
31'b0000000000000000001000000100000,
31'b0000000000000010001000000100000,
31'b0000001010110000000000000001000,
31'b0000001000000001000010000000010,
31'b0101010000000000110000000000000,
31'b0000001000100000101000000000000,
31'b0000000000100010000000100010000,
31'b0000000000100000000000100010000,
31'b1000000100000010001010000000000,
31'b1000000100000000001010000000000,
31'b0000001010100000000000000001000,
31'b0100000010000001000001100000000,
31'b0000101000000000001010001000000,
31'b0010000010100000000000100100000,
31'b0000000000000000000111000000000,
31'b0000000000110000000000100010000,
31'b0000000001100000001000000100000,
31'b1000010001000000000100000010000,
31'b0000001010010000000000000001000,
31'b0000000000001000000000100010000,
31'b0001000001000000000000100001000,
31'b0000001000000000101000000000000,
31'b0000000000000010000000100010000,
31'b0000000000000000000000100010000,
31'b0000000001010000001000000100000,
31'b0000000000000100000000100010000,
31'b0000001010000000000000000001000,
31'b0000001010000010000000000001000,
31'b0000001010000100000000000001000,
31'b0010000010000000000000100100000,
31'b0011000000000000100000000000000,
31'b0000000000010000000000100010000,
31'b0000000001000000001000000100000,
31'b0000000001000010001000000100000,
31'b1000000000000000000000011001000,
31'b1010010000000000000100000100000,
31'b1010000100000000000010100000000,
31'b1000010000000000000010010000010,
31'b1010000000000001100000000000001,
31'b0000010000000000000000010010001,
31'b0010001000100000100000100000000,
31'b0001001000110000000000000010000,
31'b0000001001100000000000000001000,
31'b0100000100000000100000001001000,
31'b0000101000001000010100000000000,
31'b0010010000000000000010000010100,
31'b0000101000000100010100000000000,
31'b0001001000100100000000000010000,
31'b0000101000000000010100000000000,
31'b0001001000100000000000000010000,
31'b0010000000000000001000000010000,
31'b0010000000000010001000000010000,
31'b0010000000000100001000000010000,
31'b0010000001010000000000100100000,
31'b0010000000001000001000000010000,
31'b0000000000000000100000000101000,
31'b0010001000000000100000100000000,
31'b0001001000010000000000000010000,
31'b0000001001000000000000000001000,
31'b0001000000000000101000100000000,
31'b0000001001000100000000000001000,
31'b0010000001000000000000100100000,
31'b0000001001001000000000000001000,
31'b0001001000000100000000000010000,
31'b0000000010000000001000000100000,
31'b0001001000000000000000000010000,
31'b0000001000110000000000000001000,
31'b0100000000010001000001100000000,
31'b0001010000000000000000010001001,
31'b0010000100000000001100000000100,
31'b0100001000000000000100100000010,
31'b0100000000000000000010010001000,
31'b1000000100000001000000001000100,
31'b1001000000000000000000011010000,
31'b0000001000100000000000000001000,
31'b0100000000000001000001100000000,
31'b0000100000000000000001000100001,
31'b0010000000100000000000100100000,
31'b0000001000101000000000000001000,
31'b0100000000010000000010010001000,
31'b0000101001000000010100000000000,
31'b0011000000000000000000001000110,
31'b0000001000010000000000000001000,
31'b0000001000010010000000000001000,
31'b0001000000000000100000000110000,
31'b0010000000010000000000100100000,
31'b0000001000011000000000000001000,
31'b0000000010000000000000100010000,
31'b0011000000000010001000000001000,
31'b0011000000000000001000000001000,
31'b0000001000000000000000000001000,
31'b0000001000000010000000000001000,
31'b0000001000000100000000000001000,
31'b0010000000000000000000100100000,
31'b0000001000001000000000000001000,
31'b0000001000001010000000000001000,
31'b0000001000001100000000000001000,
31'b0010000000001000000000100100000,
31'b0100000000000100001000001000000,
31'b0100100000010001000000000000010,
31'b0100000000000000001000001000000,
31'b0100000000000010001000001000000,
31'b0000010000000000001001000010000,
31'b1000000001000100001010000000000,
31'b0000000000000000000100100000100,
31'b1000000001000000001010000000000,
31'b0100100000000011000000000000010,
31'b0100100000000001000000000000010,
31'b0100000000010000001000001000000,
31'b0100100000000101000000000000010,
31'b1000010001100000000000000000100,
31'b0111001000000000000000001000000,
31'b0000000100100000001000000100000,
31'b1000010100000000000100000010000,
31'b0100100010000000000010000001000,
31'b1000001001000000010000000000001,
31'b0100000000100000001000001000000,
31'b0100010000000001100000000001000,
31'b1000010001010000000000000000100,
31'b1000000000000000000101000100000,
31'b0000000100010000001000000100000,
31'b1000000001100000001010000000000,
31'b1000010001001000000000000000100,
31'b1000010000000001010100000000000,
31'b0100000000000000000000000001110,
31'b0100100000000000101010000000000,
31'b1000010001000000000000000000100,
31'b1000010001000010000000000000100,
31'b0000000100000000001000000100000,
31'b0000000100000010001000000100000,
31'b0100100000000000010000000100001,
31'b0000000000000101010000100000000,
31'b0100000001000000001000001000000,
31'b0000000000000001010000100000000,
31'b1000010000110000000000000000100,
31'b1000000000000100001010000000000,
31'b1000000000000010001010000000000,
31'b1000000000000000001010000000000,
31'b1011001000000000000010000000000,
31'b0100100001000001000000000000010,
31'b0100000001010000001000001000000,
31'b0000100000000000001000010100000,
31'b1000010000100000000000000000100,
31'b1000010000100010000000000000100,
31'b1000010000100100000000000000100,
31'b1000000000010000001010000000000,
31'b1000010000011000000000000000100,
31'b1000001000000000010000000000001,
31'b0100001000000000010001000001000,
31'b0000001100000000101000000000000,
31'b1000010000010000000000000000100,
31'b0000000100000000000000100010000,
31'b1000010000010100000000000000100,
31'b1000000000100000001010000000000,
31'b1000010000001000000000000000100,
31'b1000010000001010000000000000100,
31'b1100001000000000001000010000000,
31'b0010100000000001100100000000000,
31'b1000010000000000000000000000100,
31'b1000010000000010000000000000100,
31'b1000010000000100000000000000100,
31'b1000010000000110000000000000100,
31'b1010000000000100000010100000000,
31'b1000001000000000000010000101000,
31'b1010000000000000000010100000000,
31'b1000000000000000010100001000000,
31'b0010000000000101011000000000000,
31'b0001011000000000000001000100000,
31'b0010000000000001011000000000000,
31'b1000000011000000001010000000000,
31'b0100010000100001001000000000000,
31'b0100000000000000100000001001000,
31'b1010000000010000000010100000000,
31'b1001000000000000100010000010000,
31'b1000000001000000100010000001000,
31'b0001000000000000100000000000011,
31'b0010100000000000000000110100000,
31'b0001001100100000000000000010000,
31'b0100100000000000000010000001000,
31'b0100100000000010000010000001000,
31'b1010000000100000000010100000000,
31'b1000100000000000000011000000001,
31'b0100100000001000000010000001000,
31'b0000100000000000000001000010010,
31'b0010001100000000100000100000000,
31'b0001110000000000000000000001001,
31'b0100010000000001001000000000000,
31'b0100010000000011001000000000000,
31'b0100010000000101001000000000000,
31'b1010000000000000000101000010000,
31'b1100000000000000000000010101000,
31'b0001001100000100000000000010000,
31'b0000001000000001000000010000100,
31'b0001001100000000000000000010000,
31'b0001010000010000100001000000000,
31'b0010010000000000000001100010000,
31'b1010000001000000000010100000000,
31'b0010000000000000001100000000100,
31'b1000000000010000100010000001000,
31'b1000100000100000000000001001000,
31'b1000000000000001000000001000100,
31'b1000000010000000001010000000000,
31'b0001010000000000100001000000000,
31'b0100000100000001000001100000000,
31'b0001101000000000000000010010000,
31'b0010000100100000000000100100000,
31'b1000000000000000100010000001000,
31'b1000100000000000001000000000110,
31'b1000000000010001000000001000100,
31'b1000010000000000100000001000010,
31'b0000110000000000000000000010001,
31'b1000100000001000000000001001000,
31'b0001100000000000000001000001010,
31'b0010000100010000000000100100000,
31'b1000100000000010000000001001000,
31'b1000100000000000000000001001000,
31'b1000110000000000000010000000010,
31'b1000100000000100000000001001000,
31'b0000001100000000000000000001000,
31'b0000010000000000010000101000000,
31'b0000010000000000000000010100010,
31'b0010000100000000000000100100000,
31'b1000010010000000000000000000100,
31'b1000100000010000000000001001000,
31'b1000010010000100000000000000100,
31'b0111000000000000000100000000001,
31'b1010000010000000010000000000010,
31'b0011000000100000000000000100000,
31'b0101000000000011000001000000000,
31'b0101000000000001000001000000000,
31'b1100000000000001000000001000010,
31'b0011000000101000000000000100000,
31'b0010000010100000100000100000000,
31'b1100100000010000001000000000000,
31'b0000000011100000000000000001000,
31'b0011000000110000000000000100000,
31'b0000100010001000010100000000000,
31'b1100100000001000001000000000000,
31'b0000100010000100010100000000000,
31'b1100100000000100001000000000000,
31'b0000100010000000010100000000000,
31'b1100100000000000001000000000000,
31'b0011000000000010000000000100000,
31'b0011000000000000000000000100000,
31'b0001001000000000000000100001000,
31'b0000000001000000101000000000000,
31'b0011000000001010000000000100000,
31'b0011000000001000000000000100000,
31'b0010000010000000100000100000000,
31'b0001000010010000000000000010000,
31'b0000000011000000000000000001000,
31'b0011000000010000000000000100000,
31'b0000001000001000001000000100000,
31'b0001000010001000000000000010000,
31'b0000001000000100001000000100000,
31'b0010000000000000001000100001000,
31'b0000001000000000001000000100000,
31'b0001000010000000000000000010000,
31'b0000000010110000000000000001000,
31'b0000000000000001000010000000010,
31'b0000010000000001000000001001000,
31'b0000000000100000101000000000000,
31'b0100000010000000000100100000010,
31'b0000001000100000000000100010000,
31'b1000000000000011000000000010001,
31'b1000000000000001000000000010001,
31'b0000000010100000000000000001000,
31'b0000000010100010000000000001000,
31'b0000100000000000001010001000000,
31'b0000100010000001000000000000100,
31'b0000001000000000000111000000000,
31'b0000001000110000000000100010000,
31'b0000100011000000010100000000000,
31'b1100100001000000001000000000000,
31'b0000000010010000000000000001000,
31'b0000000000000100101000000000000,
31'b0000000000000010101000000000000,
31'b0000000000000000101000000000000,
31'b0000001000000010000000100010000,
31'b0000001000000000000000100010000,
31'b0010000000000000000000000111000,
31'b0000000000001000101000000000000,
31'b0000000010000000000000000001000,
31'b0000000010000010000000000001000,
31'b0000000010000100000000000001000,
31'b0000000000010000101000000000000,
31'b0000000010001000000000000001000,
31'b0000001000010000000000100010000,
31'b0000001001000000001000000100000,
31'b0001000011000000000000000010000,
31'b1010000000000000010000000000010,
31'b1010000000000010010000000000010,
31'b1010000000000100010000000000010,
31'b0101000010000001000001000000000,
31'b1100100000000000100000000001000,
31'b0001010100000000000001000100000,
31'b0010000000100000100000100000000,
31'b0001000000110000000000000010000,
31'b0000000001100000000000000001000,
31'b0001000100000001010000000000000,
31'b0000100000001000010100000000000,
31'b0001000000101000000000000010000,
31'b0000100000000100010100000000000,
31'b0001000000100100000000000010000,
31'b0000100000000000010100000000000,
31'b0001000000100000000000000010000,
31'b0000000001010000000000000001000,
31'b0011000010000000000000000100000,
31'b0010000000001000100000100000000,
31'b0001000000011000000000000010000,
31'b0010000000000100100000100000000,
31'b0001000000010100000000000010000,
31'b0010000000000000100000100000000,
31'b0001000000010000000000000010000,
31'b0000000001000000000000000001000,
31'b0000000001000010000000000001000,
31'b0000000001000100000000000001000,
31'b0001000000001000000000000010000,
31'b0000000001001000000000000001000,
31'b0001000000000100000000000010000,
31'b0001000000000010000000000010000,
31'b0001000000000000000000000010000,
31'b0000000000110000000000000001000,
31'b0000000010000001000010000000010,
31'b0000110000000000100000000000010,
31'b0000100000010001000000000000100,
31'b0100000000000000000100100000010,
31'b0100001000000000000010010001000,
31'b0110010000000000010000000001000,
31'b1001000000000000001001000000100,
31'b0000000000100000000000000001000,
31'b0000000000100010000000000001000,
31'b0000000000100100000000000001000,
31'b0000100000000001000000000000100,
31'b0000000000101000000000000001000,
31'b0000000000101010000000000001000,
31'b0000100001000000010100000000000,
31'b0001000001100000000000000010000,
31'b0000000000010000000000000001000,
31'b0000000000010010000000000001000,
31'b0000000000010100000000000001000,
31'b0000000010000000101000000000000,
31'b0000000000011000000000000001000,
31'b0000001010000000000000100010000,
31'b0010000001000000100000100000000,
31'b0001000001010000000000000010000,
31'b0000000000000000000000000001000,
31'b0000000000000010000000000001000,
31'b0000000000000100000000000001000,
31'b0000000000000110000000000001000,
31'b0000000000001000000000000001000,
31'b0000000000001010000000000001000,
31'b0000000000001100000000000001000,
31'b0001000001000000000000000010000,
31'b0100100000001000000101000000000,
31'b1000000010000000000010000101000,
31'b0100001000000000001000001000000,
31'b0101000100000001000001000000000,
31'b0100100000000000000101000000000,
31'b0111000000010000000000001000000,
31'b0000100000000000101000010000000,
31'b1000100000000000000100000001001,
31'b1011000001000000000010000000000,
31'b0010000000000000000000000001011,
31'b1110000000000000000001000000010,
31'b0011010000000000000001000010000,
31'b0111000000000010000000001000000,
31'b0111000000000000000000001000000,
31'b0000100110000000010100000000000,
31'b1100100100000000001000000000000,
31'b1000000001000010010000000000001,
31'b1000000001000000010000000000001,
31'b0100001000100000001000001000000,
31'b0001010000000000010000001000000,
31'b1000010000000000010001000000010,
31'b1000001000000000000101000100000,
31'b0010100000000001000100000100000,
31'b0001010000001000010000001000000,
31'b1000000000000001000000000100010,
31'b1000000001010000010000000000001,
31'b1100000001000000001000010000000,
31'b0001010000010000010000001000000,
31'b1000011001000000000000000000100,
31'b0111000000100000000000001000000,
31'b0000001100000000001000000100000,
31'b0001000110000000000000000010000,
31'b1011000000010000000010000000000,
31'b1000000000100000010000000000001,
31'b0100001001000000001000001000000,
31'b0000001000000001010000100000000,
31'b0100100001000000000101000000000,
31'b1000001000000100001010000000000,
31'b1001000000000000000000010000101,
31'b1000001000000000001010000000000,
31'b1011000000000000000010000000000,
31'b1011000000000010000010000000000,
31'b1100000000100000001000010000000,
31'b0000101000000000001000010100000,
31'b0010010000000000000001000001000,
31'b0111000001000000000000001000000,
31'b0011000000000000000000000010011,
31'b1110010000000000000000000000001,
31'b1000000000000010010000000000001,
31'b1000000000000000010000000000001,
31'b0100000000000000010001000001000,
31'b0000000100000000101000000000000,
31'b1000011000010000000000000000100,
31'b1000000000001000010000000000001,
31'b0100100000000000001010000100000,
31'b0000000100001000101000000000000,
31'b0000000110000000000000000001000,
31'b1000000000010000010000000000001,
31'b1100000000000000001000010000000,
31'b0000000100010000101000000000000,
31'b1000011000000000000000000000100,
31'b1000011000000010000000000000100,
31'b1100000000001000001000010000000,
31'b0001000111000000000000000010000,
31'b1010000100000000010000000000010,
31'b1000000000000000000010000101000,
31'b1010001000000000000010100000000,
31'b1000001000000000010100001000000,
31'b0100100010000000000101000000000,
31'b0001010000000000000001000100000,
31'b0010001000000001011000000000000,
31'b0001010000000100000001000100000,
31'b0001000000000011010000000000000,
31'b0001000000000001010000000000000,
31'b0001100001000000000000010010000,
31'b0001000000000101010000000000000,
31'b0001000001000000000100000000100,
31'b0000100000000000000000010001000,
31'b0000100100000000010100000000000,
31'b0001000100100000000000000010000,
31'b0010000000000001000010000000001,
31'b1000000011000000010000000000001,
31'b0010000100001000100000100000000,
31'b0001010010000000010000001000000,
31'b0010000100000100100000100000000,
31'b0001010000100000000001000100000,
31'b0010000100000000100000100000000,
31'b0001000100010000000000000010000,
31'b0000000101000000000000000001000,
31'b0001000000100001010000000000000,
31'b0000000101000100000000000001000,
31'b0001000100001000000000000010000,
31'b0000000101001000000000000001000,
31'b0001000100000100000000000010000,
31'b0000000000000001000000010000100,
31'b0001000100000000000000000010000,
31'b0001000000000000000000000100011,
31'b1000000010100000010000000000001,
31'b0001100000010000000000010010000,
31'b0010100000000000100000110000000,
31'b0100000000000000000000001101000,
31'b0110010000000000000100010000000,
31'b1001000000000000000010000110000,
31'b1000001010000000001010000000000,
31'b0000000100100000000000000001000,
31'b0001000001000001010000000000000,
31'b0001100000000000000000010010000,
31'b0000100100000001000000000000100,
31'b0001000000000000000100000000100,
31'b0001000000000010000100000000100,
31'b0001000000000100000100000000100,
31'b0001000101100000000000000010000,
31'b0000000100010000000000000001000,
31'b1000000010000000010000000000001,
31'b0000000100010100000000000001000,
31'b0000000110000000101000000000000,
31'b0000000100011000000000000001000,
31'b1000101000000000000000001001000,
31'b0010000101000000100000100000000,
31'b0001010000000000001110000000000,
31'b0000000100000000000000000001000,
31'b0000000100000010000000000001000,
31'b0000000100000100000000000001000,
31'b0000000000000000010100010000000,
31'b0000000100001000000000000001000,
31'b0000100000000000010000000010100,
31'b0000000100001100000000000001000,
31'b0001000101000000000000000010000,
31'b0110000000000000011000000100000,
31'b0010100000000000000000000010010,
31'b0101000001000000110000000000000,
31'b1000000010000000000010010000010,
31'b0000000100000000001001000010000,
31'b0000000000000000000010000100100,
31'b1000000000100000000011100000000,
31'b1000000000010000000100000010000,
31'b1001000001000000000100000001000,
31'b1000100000000000000000010000100,
31'b1000000000100001000000010001000,
31'b1000000000001000000100000010000,
31'b1000000101100000000000000000100,
31'b1000000000000100000100000010000,
31'b1000000000000010000100000010000,
31'b1000000000000000000100000010000,
31'b0011000000000000010100000000010,
31'b0011011000000000000000000100000,
31'b0001010000000000000000100001000,
31'b0100000100000001100000000001000,
31'b1000000101010000000000000000100,
31'b0000010001000000000000100010000,
31'b1000000000000000000011100000000,
31'b1000000000110000000100000010000,
31'b1000000101001000000000000000100,
31'b1000100000100000000000010000100,
31'b1000000000000001000000010001000,
31'b1000000000101000000100000010000,
31'b1000000101000000000000000000100,
31'b1000000101000010000000000000100,
31'b0000010000000000001000000100000,
31'b1000000000100000000100000010000,
31'b1100000000000000000000001100100,
31'b0010100001000000000000000010010,
31'b0101000000000000110000000000000,
31'b0101000000000010110000000000000,
31'b1000000100110000000000000000100,
31'b0000010000100000000000100010000,
31'b0101000000001000110000000000000,
31'b1000010100000000001010000000000,
31'b1001000000000000000100000001000,
31'b1001000000000010000100000001000,
31'b1001000000000100000100000001000,
31'b1001000100000000010000010000000,
31'b1000000100100000000000000000100,
31'b1000000100100010000000000000100,
31'b1000000100100100000000000000100,
31'b1000000001000000000100000010000,
31'b1000000100011000000000000000100,
31'b0000101000000000000000001000100,
31'b0101000000100000110000000000000,
31'b0100000000000000000001101000000,
31'b1000000100010000000000000000100,
31'b0000010000000000000000100010000,
31'b1000000100010100000000000000100,
31'b0000010000000100000000100010000,
31'b1000000100001000000000000000100,
31'b1000100000000000010000000011000,
31'b1000000100001100000000000000100,
31'b0110000000000000100010000000001,
31'b1000000100000000000000000000100,
31'b1000000100000010000000000000100,
31'b1000000100000100000000000000100,
31'b1000000100000110000000000000100,
31'b1010000000000010000100000100000,
31'b1010000000000000000100000100000,
31'b1000001000000000000100100001000,
31'b1000000000000000000010010000010,
31'b0000000000000010000000010010001,
31'b0000000000000000000000010010001,
31'b0100000001000000000000011000010,
31'b0000100000010000000000000100010,
31'b0100001000000000110000100000000,
31'b1010000000010000000100000100000,
31'b0100000100000000100010000000010,
31'b0010000000000000000010000010100,
31'b0100000000000100011000000010000,
31'b0000100000000100000000000100010,
31'b0100000000000000011000000010000,
31'b0000100000000000000000000100010,
31'b0010010000000000001000000010000,
31'b1010000000100000000100000100000,
31'b0010010000000100001000000010000,
31'b1100000000000001000101000000000,
31'b0010010000001000001000000010000,
31'b0000010000000000100000000101000,
31'b1100001000010000000000000000010,
31'b0001100100000000000000000001001,
31'b0100000100000001001000000000000,
31'b0101001000000000000001001000000,
31'b1100001000001000000000000000010,
31'b0010010001000000000000100100000,
31'b1100001000000100000000000000010,
31'b0001100000000000100001010000000,
31'b1100001000000000000000000000010,
31'b0001011000000000000000000010000,
31'b0001000100010000100001000000000,
31'b1101000000000000000001010000000,
31'b0001000000000000000000010001001,
31'b1001000000000000101100000000000,
31'b0100000000000100000000011000010,
31'b0100000000000000010000100100000,
31'b0100000000000000000000011000010,
31'b0100000000000100010000100100000,
31'b0001000100000000100001000000000,
31'b0101000000000000011000000001000,
31'b0001000100000100100001000000000,
31'b0010010000100000000000100100000,
31'b1010001000000000100100000000000,
31'b0100100000000001001000010000000,
31'b0100000001000000011000000010000,
31'b0000100001000000000000000100010,
31'b0000100100000000000000000010001,
31'b0000101010000000000000001000100,
31'b0001010000000000100000000110000,
31'b1100000000000000100000000100010,
31'b1000101000000000010000100000000,
31'b0000010010000000000000100010000,
31'b1100000000000000010001000000100,
31'b0011010000000000001000000001000,
31'b0000011000000000000000000001000,
31'b0000011000000010000000000001000,
31'b0000011000000100000000000001000,
31'b0010010000000000000000100100000,
31'b1000000110000000000000000000100,
31'b1000001000000000000000001010001,
31'b1100001001000000000000000000010,
31'b0011100000000001000010000000000,
31'b0100100000000000100000000000100,
31'b0100100000000010100000000000100,
31'b0100010000000000001000001000000,
31'b0100010000000010001000001000000,
31'b0000000000000000001001000010000,
31'b0000000100000000000010000100100,
31'b0000010000000000000100100000100,
31'b1000010001000000001010000000000,
31'b1001100000000001000000000010000,
31'b1000100100000000000000010000100,
31'b0100010000010000001000001000000,
31'b1001000001000000010000010000000,
31'b1000000001100000000000000000100,
31'b1000000100000100000100000010000,
31'b1000000100000010000100000010000,
31'b1000000100000000000100000010000,
31'b1000000001011000000000000000100,
31'b1000001000000000100000000100100,
31'b0100010000100000001000001000000,
31'b0100000000000001100000000001000,
31'b1000000001010000000000000000100,
31'b1000010000000000000101000100000,
31'b1000000100000000000011100000000,
31'b0110000000000000000000011000001,
31'b1000000001001000000000000000100,
31'b1000000000000001010100000000000,
31'b1000000100000001000000010001000,
31'b1001000000000000000000000011100,
31'b1000000001000000000000000000100,
31'b1000000001000010000000000000100,
31'b1000000001000100000000000000100,
31'b1000000100100000000100000010000,
31'b1101000000000000001000000000001,
31'b0010000010000000000001100010000,
31'b0101000100000000110000000000000,
31'b0001000000000000001001000001000,
31'b1000000000110000000000000000100,
31'b1000010000000100001010000000000,
31'b1000010000000010001010000000000,
31'b1000010000000000001010000000000,
31'b1000000000101000000000000000100,
31'b1001000000000100010000010000000,
31'b1001000000000010010000010000000,
31'b1001000000000000010000010000000,
31'b1000000000100000000000000000100,
31'b1000000000100010000000000000100,
31'b1000000000100100000000000000100,
31'b0000000000000000000001100100000,
31'b1000000000011000000000000000100,
31'b1000011000000000010000000000001,
31'b1010000000000000000010010000001,
31'b0100000100000000000001101000000,
31'b1000000000010000000000000000100,
31'b1000000000010010000000000000100,
31'b1000000000010100000000000000100,
31'b1000010000100000001010000000000,
31'b1000000000001000000000000000100,
31'b1000000000001010000000000000100,
31'b1000000000001100000000000000100,
31'b1001000000100000010000010000000,
31'b1000000000000000000000000000100,
31'b1000000000000010000000000000100,
31'b1000000000000100000000000000100,
31'b1000000000000110000000000000100,
31'b0100100010000000100000000000100,
31'b1010000100000000000100000100000,
31'b1010010000000000000010100000000,
31'b1000010000000000010100001000000,
31'b0001000000000001000000000000101,
31'b0001001000000000000001000100000,
31'b0011000000000000000001100001000,
31'b0001100000100000000000000001001,
31'b0100000000100001001000000000000,
31'b0100010000000000100000001001000,
31'b0100000000000000100010000000010,
31'b0100100000000000001000000001100,
31'b1100000000000000100000000010001,
31'b0001010000000000100000000000011,
31'b0100000100000000011000000010000,
31'b0000100100000000000000000100010,
31'b0100000000010001001000000000000,
31'b0100100000000100000000001000010,
31'b0100100000000010000000001000010,
31'b0100100000000000000000001000010,
31'b1101100000000000000001000000000,
31'b0001100000000100000000000001001,
31'b1001001000000000000000100000100,
31'b0001100000000000000000000001001,
31'b0100000000000001001000000000000,
31'b0100000000000011001000000000000,
31'b0100000000000101001000000000000,
31'b0100100000010000000000001000010,
31'b1000000011000000000000000000100,
31'b1110000000000000000100001000000,
31'b1100001100000000000000000000010,
31'b0001100000010000000000000001001,
31'b0001000000010000100001000000000,
31'b0010000000000000000001100010000,
31'b0001000100000000000000010001001,
31'b0010010000000000001100000000100,
31'b1000100000000001101000000000000,
31'b0110001000000000000100010000000,
31'b1000100000100000000010000000010,
31'b1000010010000000001010000000000,
31'b0001000000000000100001000000000,
31'b0001000000000010100001000000000,
31'b0001000000000100100001000000000,
31'b1001000010000000010000010000000,
31'b1000000010100000000000000000100,
31'b1000000010100010000000000000100,
31'b1000000010100100000000000000100,
31'b1000000000000000100000001000010,
31'b0000100000000000000000000010001,
31'b0000100000000010000000000010001,
31'b0000100000000100000000000010001,
31'b0100100001000000000000001000010,
31'b1000000010010000000000000000100,
31'b1000110000000000000000001001000,
31'b1000100000000000000010000000010,
31'b1000100000000010000010000000010,
31'b0010000000000000000110000000000,
31'b0000000000000000010000101000000,
31'b0000000000000000000000010100010,
31'b0000000000000100010000101000000,
31'b1000000010000000000000000000100,
31'b1000000010000010000000000000100,
31'b1000000010000100000000000000100,
31'b1000000010000110000000000000100,
31'b0000000100001000000000011000100,
31'b0011010000100000000000000100000,
31'b0000000100000000100001100000000,
31'b0101010000000001000001000000000,
31'b0000000100000000000000011000100,
31'b0001000000000001000000001010000,
31'b0010000001000000100000010000001,
31'b1100000000000001000010000001000,
31'b0000000001000000100010000000100,
31'b1000101000000000000000010000100,
31'b0010000100000000000010001000001,
31'b1100000000000000000001110000000,
31'b0010000101000000000001000001000,
31'b1100000000000000100000001000100,
31'b1100000010100000000000000000010,
31'b1000001000000000000100000010000,
31'b0110100010000000000100000000000,
31'b0011010000000000000000000100000,
31'b0001011000000000000000100001000,
31'b0001000100000000010000001000000,
31'b1100100000000000000010000000100,
31'b0011010000001000000000000100000,
31'b1100000010010000000000000000010,
31'b0001010010010000000000000010000,
31'b0100000000000000000000010100100,
31'b0101000010000000000001001000000,
31'b1100000010001000000000000000010,
31'b0001010010001000000000000010000,
31'b1100000010000100000000000000010,
31'b0011000000000001010001000000000,
31'b1100000010000000000000000000010,
31'b0001010010000000000000000010000,
31'b0000000000010000100010000000100,
31'b0000100000100000000000001000100,
31'b0000000000000001000000001001000,
31'b0000010000100000101000000000000,
31'b0010000100010000000001000001000,
31'b0001100000000000000000100100010,
31'b0010000000000000100000010000001,
31'b1010000000000000001100000001000,
31'b0000000000000000100010000000100,
31'b0000100000000000001000000001010,
31'b0000000000010001000000001001000,
31'b0000110010000001000000000000100,
31'b0010000100000000000001000001000,
31'b0110000000000000111000000000000,
31'b0010000100000100000001000001000,
31'b1110000100000000000000000000001,
31'b0000100000000010000000001000100,
31'b0000100000000000000000001000100,
31'b0000010000000010101000000000000,
31'b0000010000000000101000000000000,
31'b1000100010000000010000100000000,
31'b0000100000001000000000001000100,
31'b0010010000000000000000000111000,
31'b0000010000001000101000000000000,
31'b0000010010000000000000000001000,
31'b0000100000010000000000001000100,
31'b0000010010000100000000000001000,
31'b0000010000010000101000000000000,
31'b1000001100000000000000000000100,
31'b1000001100000010000000000000100,
31'b1100000011000000000000000000010,
31'b0001010011000000000000000010000,
31'b1010010000000000010000000000010,
31'b1010001000000000000100000100000,
31'b1000000000000000000100100001000,
31'b1000001000000000000010010000010,
31'b0001000100000010000001000100000,
31'b0001000100000000000001000100000,
31'b1100000000110000000000000000010,
31'b0001010000110000000000000010000,
31'b0100000000000000110000100000000,
31'b0101000000100000000001001000000,
31'b1100000000101000000000000000010,
31'b0011000000000001000000001100000,
31'b1100000000100100000000000000010,
31'b0001010000100100000000000010000,
31'b1100000000100000000000000000010,
31'b0001010000100000000000000010000,
31'b0110100000000000000100000000000,
31'b0110100000000010000100000000000,
31'b1100000000011000000000000000010,
31'b0001010000011000000000000010000,
31'b1100000000010100000000000000010,
31'b0001010000010100000000000010000,
31'b1100000000010000000000000000010,
31'b0001010000010000000000000010000,
31'b0000010001000000000000000001000,
31'b0101000000000000000001001000000,
31'b1100000000001000000000000000010,
31'b0001010000001000000000000010000,
31'b1100000000000100000000000000010,
31'b0001010000000100000000000010000,
31'b1100000000000000000000000000010,
31'b0001010000000000000000000010000,
31'b0000100000000100100000000000010,
31'b0000100010100000000000001000100,
31'b0000100000000000100000000000010,
31'b0000100000000010100000000000010,
31'b1010000000010000100100000000000,
31'b1010000000000000010001000000001,
31'b0110000000000000010000000001000,
31'b0110000000000010010000000001000,
31'b0000010000100000000000000001000,
31'b0000010000100010000000000001000,
31'b0000100000010000100000000000010,
31'b0000110000000001000000000000100,
31'b1010000000000000100100000000000,
31'b1010000000000010100100000000000,
31'b1100000001100000000000000000010,
31'b0001010001100000000000000010000,
31'b0000010000010000000000000001000,
31'b0000100010000000000000001000100,
31'b0000100000100000100000000000010,
31'b0000010010000000101000000000000,
31'b1000100000000000010000100000000,
31'b1000100000000010010000100000000,
31'b1100000001010000000000000000010,
31'b0001010001010000000000000010000,
31'b0000010000000000000000000001000,
31'b0000010000000010000000000001000,
31'b0000010000000100000000000001000,
31'b0000000000000000000010001000010,
31'b0000010000001000000000000001000,
31'b1000000000000000000000001010001,
31'b1100000001000000000000000000010,
31'b0001010001000000000000000010000,
31'b0000000000001000000000011000100,
31'b1000000010000000010000110000000,
31'b0000000000000000100001100000000,
31'b0001000000100000010000001000000,
31'b0000000000000000000000011000100,
31'b0001000010000000000001000100000,
31'b0000000000001000100001100000000,
31'b0001000010000100000001000100000,
31'b0010000001001000000001000001000,
31'b0011000000000100000001000010000,
31'b0010000000000000000010001000001,
31'b0011000000000000000001000010000,
31'b0010000001000000000001000001000,
31'b0111010000000000000000001000000,
31'b0010000001000100000001000001000,
31'b1110000001000000000000000000001,
31'b1000000000001000010001000000010,
31'b1000000000000000100000000100100,
31'b0001000000000010010000001000000,
31'b0001000000000000010000001000000,
31'b1000000000000000010001000000010,
31'b1000000000001000100000000100100,
31'b1001000010000000000000100000100,
31'b0001000000001000010000001000000,
31'b1000010000000001000000000100010,
31'b1000001000000001010100000000000,
31'b0010100000000000010101000000000,
31'b0001000000010000010000001000000,
31'b1000001001000000000000000000100,
31'b1000001001000010000000000000100,
31'b1100000110000000000000000000010,
31'b0001010110000000000000000010000,
31'b0010000000011000000001000001000,
31'b1100000000000000000010010000100,
31'b0000000100000001000000001001000,
31'b0001001000000000001001000001000,
31'b0010000000010000000001000001000,
31'b0110000010000000000100010000000,
31'b0010000100000000100000010000001,
31'b1110000000010000000000000000001,
31'b0010000000001000000001000001000,
31'b0110000000000000000010000010010,
31'b0010000001000000000010001000001,
31'b1110000000001000000000000000001,
31'b0010000000000000000001000001000,
31'b0100100000000000000000000100100,
31'b0010000000000100000001000001000,
31'b1110000000000000000000000000001,
31'b1000010000000010010000000000001,
31'b1000010000000000010000000000001,
31'b0101000000000001001000100000000,
31'b0001000001000000010000001000000,
31'b1000001000010000000000000000100,
31'b1000010000001000010000000000001,
31'b1101000000000000010010000000000,
31'b0001000010000000001110000000000,
31'b1000001000001000000000000000100,
31'b1000010000010000010000000000001,
31'b1100010000000000001000010000000,
31'b0001000001010000010000001000000,
31'b1000001000000000000000000000100,
31'b1000001000000010000000000000100,
31'b1000001000000100000000000000100,
31'b1110000000100000000000000000001,
31'b1000000000000100000000001100010,
31'b1000000000000000010000110000000,
31'b1000000000000000000000001100010,
31'b1000000000000100010000110000000,
31'b0001000000000010000001000100000,
31'b0001000000000000000001000100000,
31'b1001000000100000000000100000100,
31'b0001000000000100000001000100000,
31'b0100001000100001001000000000000,
31'b0001010000000001010000000000000,
31'b1100000000000000001000100000001,
31'b0011000010000000000001000010000,
31'b0010100000000000000100001100000,
31'b0001000000010000000001000100000,
31'b1100000100100000000000000000010,
31'b0001010100100000000000000010000,
31'b0110100100000000000100000000000,
31'b1000000010000000100000000100100,
31'b1001000000001000000000100000100,
31'b0001000010000000010000001000000,
31'b1001000000000100000000100000100,
31'b0001000000100000000001000100000,
31'b1001000000000000000000100000100,
31'b0000000000000000100000010000010,
31'b0100001000000001001000000000000,
31'b0101000100000000000001001000000,
31'b1100000100001000000000000000010,
31'b0001010100001000000000000010000,
31'b1100000100000100000000000000010,
31'b0001010100000100000000000010000,
31'b1100000100000000000000000000010,
31'b0001010100000000000000000010000,
31'b0001010000000000000000000100011,
31'b1100000000000000000000000110001,
31'b0000100100000000100000000000010,
31'b0110100000000000000000000010100,
31'b0110000000000010000100010000000,
31'b0110000000000000000100010000000,
31'b0110000100000000010000000001000,
31'b0100000000000000000010000100010,
31'b0001001000000000100001000000000,
31'b0001010001000001010000000000000,
31'b0001110000000000000000010010000,
31'b1100100000000000000000010000010,
31'b0010000010000000000001000001000,
31'b0110000000010000000100010000000,
31'b0010000010000100000001000001000,
31'b1110000010000000000000000000001,
31'b0000101000000000000000000010001,
31'b1000010010000000010000000000001,
31'b0000101000000100000000000010001,
31'b0001000011000000010000001000000,
31'b1000100100000000010000100000000,
31'b0110000000100000000100010000000,
31'b1001000001000000000000100000100,
31'b0001000000000000001110000000000,
31'b0000010100000000000000000001000,
31'b0000010100000010000000000001000,
31'b0000010100000100000000000001000,
31'b0000010000000000010100010000000,
31'b1000001010000000000000000000100,
31'b1000001010000010000000000000100,
31'b1100000101000000000000000000010,
31'b0001010101000000000000000010000
};

